magic
tech sky130A
magscale 1 2
timestamp 1743983958
<< checkpaint >>
rect -3932 -3932 27400 29544
<< viali >>
rect 7389 23273 7423 23307
rect 8033 23273 8067 23307
rect 11621 23273 11655 23307
rect 14473 23273 14507 23307
rect 17417 23273 17451 23307
rect 18337 23273 18371 23307
rect 9321 23205 9355 23239
rect 12265 23205 12299 23239
rect 16957 23205 16991 23239
rect 18797 23205 18831 23239
rect 13185 23137 13219 23171
rect 16221 23137 16255 23171
rect 4813 23069 4847 23103
rect 5273 23069 5307 23103
rect 6561 23069 6595 23103
rect 8677 23069 8711 23103
rect 9137 23069 9171 23103
rect 9781 23069 9815 23103
rect 10425 23069 10459 23103
rect 11069 23069 11103 23103
rect 13461 23069 13495 23103
rect 13737 23069 13771 23103
rect 15117 23069 15151 23103
rect 15577 23069 15611 23103
rect 16037 23069 16071 23103
rect 17969 23069 18003 23103
rect 18981 23069 19015 23103
rect 19441 23069 19475 23103
rect 7297 23001 7331 23035
rect 7941 23001 7975 23035
rect 11897 23001 11931 23035
rect 12449 23001 12483 23035
rect 13001 23001 13035 23035
rect 14381 23001 14415 23035
rect 16773 23001 16807 23035
rect 17325 23001 17359 23035
rect 18245 23001 18279 23035
rect 4629 22933 4663 22967
rect 5457 22933 5491 22967
rect 6745 22933 6779 22967
rect 8493 22933 8527 22967
rect 9965 22933 9999 22967
rect 10609 22933 10643 22967
rect 11253 22933 11287 22967
rect 12633 22933 12667 22967
rect 13093 22933 13127 22967
rect 13645 22933 13679 22967
rect 13921 22933 13955 22967
rect 14933 22933 14967 22967
rect 15393 22933 15427 22967
rect 15669 22933 15703 22967
rect 16129 22933 16163 22967
rect 17785 22933 17819 22967
rect 19625 22933 19659 22967
rect 7757 22729 7791 22763
rect 13599 22729 13633 22763
rect 15347 22729 15381 22763
rect 7849 22661 7883 22695
rect 8539 22661 8573 22695
rect 13185 22661 13219 22695
rect 15853 22661 15887 22695
rect 1501 22593 1535 22627
rect 8366 22593 8400 22627
rect 8642 22593 8676 22627
rect 13093 22593 13127 22627
rect 13670 22593 13704 22627
rect 15276 22593 15310 22627
rect 15945 22593 15979 22627
rect 16359 22593 16393 22627
rect 16462 22593 16496 22627
rect 16681 22593 16715 22627
rect 2053 22525 2087 22559
rect 8033 22525 8067 22559
rect 13369 22525 13403 22559
rect 16083 22525 16117 22559
rect 7389 22389 7423 22423
rect 8263 22389 8297 22423
rect 12725 22389 12759 22423
rect 15485 22389 15519 22423
rect 16865 22389 16899 22423
rect 13553 22117 13587 22151
rect 7941 22049 7975 22083
rect 8585 22049 8619 22083
rect 13277 22049 13311 22083
rect 14151 22049 14185 22083
rect 14749 22049 14783 22083
rect 14933 22049 14967 22083
rect 15577 22049 15611 22083
rect 15853 22049 15887 22083
rect 16129 22049 16163 22083
rect 1409 21981 1443 22015
rect 6929 21981 6963 22015
rect 7297 21981 7331 22015
rect 7849 21981 7883 22015
rect 8401 21981 8435 22015
rect 12265 21981 12299 22015
rect 13185 21981 13219 22015
rect 13737 21981 13771 22015
rect 14238 21981 14272 22015
rect 16221 21981 16255 22015
rect 7113 21913 7147 21947
rect 7757 21913 7791 21947
rect 8217 21913 8251 21947
rect 12449 21913 12483 21947
rect 12633 21913 12667 21947
rect 13093 21913 13127 21947
rect 13921 21913 13955 21947
rect 14565 21913 14599 21947
rect 15393 21913 15427 21947
rect 1593 21845 1627 21879
rect 7389 21845 7423 21879
rect 12725 21845 12759 21879
rect 15025 21845 15059 21879
rect 15485 21845 15519 21879
rect 5181 21641 5215 21675
rect 8033 21641 8067 21675
rect 15945 21641 15979 21675
rect 16313 21573 16347 21607
rect 1501 21505 1535 21539
rect 4502 21505 4536 21539
rect 5273 21505 5307 21539
rect 5687 21505 5721 21539
rect 5790 21505 5824 21539
rect 7113 21505 7147 21539
rect 7941 21505 7975 21539
rect 8585 21505 8619 21539
rect 12817 21505 12851 21539
rect 15669 21505 15703 21539
rect 16129 21505 16163 21539
rect 5457 21437 5491 21471
rect 7205 21437 7239 21471
rect 8125 21437 8159 21471
rect 12725 21437 12759 21471
rect 13461 21437 13495 21471
rect 15485 21437 15519 21471
rect 1685 21369 1719 21403
rect 8401 21369 8435 21403
rect 13277 21369 13311 21403
rect 4399 21301 4433 21335
rect 4813 21301 4847 21335
rect 7481 21301 7515 21335
rect 7573 21301 7607 21335
rect 8769 21301 8803 21335
rect 13185 21301 13219 21335
rect 13645 21301 13679 21335
rect 15853 21301 15887 21335
rect 15209 21029 15243 21063
rect 4537 20961 4571 20995
rect 4721 20961 4755 20995
rect 7297 20961 7331 20995
rect 18613 20961 18647 20995
rect 19901 20961 19935 20995
rect 1685 20893 1719 20927
rect 4905 20893 4939 20927
rect 7481 20893 7515 20927
rect 8309 20893 8343 20927
rect 13461 20893 13495 20927
rect 13829 20893 13863 20927
rect 15393 20893 15427 20927
rect 15577 20893 15611 20927
rect 16129 20893 16163 20927
rect 16313 20893 16347 20927
rect 17417 20893 17451 20927
rect 17509 20893 17543 20927
rect 18429 20893 18463 20927
rect 18889 20893 18923 20927
rect 19625 20893 19659 20927
rect 20202 20893 20236 20927
rect 22017 20893 22051 20927
rect 4445 20825 4479 20859
rect 5181 20825 5215 20859
rect 5641 20825 5675 20859
rect 5825 20825 5859 20859
rect 7665 20825 7699 20859
rect 8125 20825 8159 20859
rect 13645 20825 13679 20859
rect 15945 20825 15979 20859
rect 17969 20825 18003 20859
rect 19073 20825 19107 20859
rect 1501 20757 1535 20791
rect 4077 20757 4111 20791
rect 5457 20757 5491 20791
rect 7941 20757 7975 20791
rect 18245 20757 18279 20791
rect 18705 20757 18739 20791
rect 19257 20757 19291 20791
rect 19717 20757 19751 20791
rect 20131 20757 20165 20791
rect 21833 20757 21867 20791
rect 5273 20553 5307 20587
rect 10793 20553 10827 20587
rect 18337 20553 18371 20587
rect 18429 20553 18463 20587
rect 19257 20553 19291 20587
rect 4261 20485 4295 20519
rect 5825 20485 5859 20519
rect 13645 20485 13679 20519
rect 19625 20485 19659 20519
rect 4537 20417 4571 20451
rect 5365 20417 5399 20451
rect 6009 20417 6043 20451
rect 6193 20417 6227 20451
rect 7297 20417 7331 20451
rect 9321 20417 9355 20451
rect 9413 20417 9447 20451
rect 10885 20417 10919 20451
rect 11575 20417 11609 20451
rect 11662 20417 11696 20451
rect 13185 20417 13219 20451
rect 15301 20417 15335 20451
rect 17141 20417 17175 20451
rect 18981 20417 19015 20451
rect 19717 20417 19751 20451
rect 20131 20417 20165 20451
rect 20234 20417 20268 20451
rect 3893 20349 3927 20383
rect 4077 20349 4111 20383
rect 4629 20349 4663 20383
rect 5181 20349 5215 20383
rect 7205 20349 7239 20383
rect 9873 20349 9907 20383
rect 10977 20349 11011 20383
rect 13093 20349 13127 20383
rect 15393 20349 15427 20383
rect 17233 20349 17267 20383
rect 18521 20349 18555 20383
rect 19901 20349 19935 20383
rect 19165 20281 19199 20315
rect 4905 20213 4939 20247
rect 5733 20213 5767 20247
rect 7665 20213 7699 20247
rect 10425 20213 10459 20247
rect 14933 20213 14967 20247
rect 16773 20213 16807 20247
rect 17969 20213 18003 20247
rect 18797 20213 18831 20247
rect 5273 20009 5307 20043
rect 15853 20009 15887 20043
rect 17877 20009 17911 20043
rect 10701 19941 10735 19975
rect 12817 19941 12851 19975
rect 5641 19873 5675 19907
rect 6009 19873 6043 19907
rect 7849 19873 7883 19907
rect 8953 19873 8987 19907
rect 9413 19873 9447 19907
rect 9689 19873 9723 19907
rect 10149 19873 10183 19907
rect 11345 19873 11379 19907
rect 12265 19873 12299 19907
rect 13461 19873 13495 19907
rect 15485 19873 15519 19907
rect 16589 19873 16623 19907
rect 17233 19873 17267 19907
rect 18337 19873 18371 19907
rect 1685 19805 1719 19839
rect 4997 19805 5031 19839
rect 5089 19805 5123 19839
rect 5825 19805 5859 19839
rect 7573 19805 7607 19839
rect 7665 19805 7699 19839
rect 8033 19805 8067 19839
rect 9321 19805 9355 19839
rect 10057 19805 10091 19839
rect 12449 19805 12483 19839
rect 13369 19805 13403 19839
rect 13737 19805 13771 19839
rect 14657 19805 14691 19839
rect 15209 19805 15243 19839
rect 15301 19805 15335 19839
rect 16037 19805 16071 19839
rect 16773 19805 16807 19839
rect 18245 19805 18279 19839
rect 18705 19805 18739 19839
rect 18889 19805 18923 19839
rect 22017 19805 22051 19839
rect 11529 19737 11563 19771
rect 11713 19737 11747 19771
rect 12357 19737 12391 19771
rect 14473 19737 14507 19771
rect 15761 19737 15795 19771
rect 16681 19737 16715 19771
rect 1501 19669 1535 19703
rect 7205 19669 7239 19703
rect 11069 19669 11103 19703
rect 11161 19669 11195 19703
rect 11897 19669 11931 19703
rect 12909 19669 12943 19703
rect 13277 19669 13311 19703
rect 14841 19669 14875 19703
rect 17141 19669 17175 19703
rect 18521 19669 18555 19703
rect 21833 19669 21867 19703
rect 7297 19465 7331 19499
rect 7389 19465 7423 19499
rect 8769 19465 8803 19499
rect 10149 19465 10183 19499
rect 10241 19465 10275 19499
rect 11575 19465 11609 19499
rect 13553 19465 13587 19499
rect 14013 19465 14047 19499
rect 14289 19465 14323 19499
rect 14657 19465 14691 19499
rect 14749 19465 14783 19499
rect 16681 19465 16715 19499
rect 17049 19465 17083 19499
rect 17141 19465 17175 19499
rect 21833 19465 21867 19499
rect 9321 19397 9355 19431
rect 10609 19397 10643 19431
rect 10793 19397 10827 19431
rect 1685 19329 1719 19363
rect 5181 19329 5215 19363
rect 11646 19329 11680 19363
rect 13093 19329 13127 19363
rect 13737 19329 13771 19363
rect 13829 19329 13863 19363
rect 22017 19329 22051 19363
rect 5089 19261 5123 19295
rect 7205 19261 7239 19295
rect 8309 19261 8343 19295
rect 8861 19261 8895 19295
rect 9045 19261 9079 19295
rect 9505 19261 9539 19295
rect 9689 19261 9723 19295
rect 10333 19261 10367 19295
rect 13185 19261 13219 19295
rect 13461 19261 13495 19295
rect 14933 19261 14967 19295
rect 17325 19261 17359 19295
rect 1501 19125 1535 19159
rect 5549 19125 5583 19159
rect 7757 19125 7791 19159
rect 8401 19125 8435 19159
rect 9781 19125 9815 19159
rect 10977 19125 11011 19159
rect 5089 18921 5123 18955
rect 6469 18921 6503 18955
rect 10057 18921 10091 18955
rect 2881 18785 2915 18819
rect 4261 18785 4295 18819
rect 6193 18785 6227 18819
rect 8401 18785 8435 18819
rect 8585 18785 8619 18819
rect 10425 18785 10459 18819
rect 1409 18717 1443 18751
rect 2421 18717 2455 18751
rect 2605 18717 2639 18751
rect 3065 18717 3099 18751
rect 4445 18717 4479 18751
rect 5181 18717 5215 18751
rect 5917 18717 5951 18751
rect 6009 18717 6043 18751
rect 6745 18717 6779 18751
rect 8309 18717 8343 18751
rect 10241 18717 10275 18751
rect 18153 18717 18187 18751
rect 22017 18717 22051 18751
rect 3249 18649 3283 18683
rect 4721 18649 4755 18683
rect 4905 18649 4939 18683
rect 6561 18649 6595 18683
rect 1593 18581 1627 18615
rect 2789 18581 2823 18615
rect 4629 18581 4663 18615
rect 5549 18581 5583 18615
rect 7941 18581 7975 18615
rect 21833 18581 21867 18615
rect 2513 18377 2547 18411
rect 3249 18377 3283 18411
rect 3341 18377 3375 18411
rect 5641 18377 5675 18411
rect 5733 18377 5767 18411
rect 7205 18377 7239 18411
rect 7757 18377 7791 18411
rect 13553 18377 13587 18411
rect 16037 18377 16071 18411
rect 17325 18377 17359 18411
rect 17693 18377 17727 18411
rect 18153 18377 18187 18411
rect 18705 18377 18739 18411
rect 19993 18377 20027 18411
rect 4353 18309 4387 18343
rect 14013 18309 14047 18343
rect 17233 18309 17267 18343
rect 19073 18309 19107 18343
rect 19717 18309 19751 18343
rect 19901 18309 19935 18343
rect 20361 18309 20395 18343
rect 1685 18241 1719 18275
rect 1904 18241 1938 18275
rect 3893 18241 3927 18275
rect 4905 18241 4939 18275
rect 7389 18241 7423 18275
rect 7573 18241 7607 18275
rect 13093 18241 13127 18275
rect 13185 18241 13219 18275
rect 13369 18241 13403 18275
rect 13645 18241 13679 18275
rect 13921 18241 13955 18275
rect 15853 18241 15887 18275
rect 16129 18241 16163 18275
rect 18061 18241 18095 18275
rect 19165 18241 19199 18275
rect 19533 18241 19567 18275
rect 20453 18241 20487 18275
rect 20867 18241 20901 18275
rect 20970 18241 21004 18275
rect 21373 18241 21407 18275
rect 2329 18173 2363 18207
rect 2421 18173 2455 18207
rect 3157 18173 3191 18207
rect 3801 18173 3835 18207
rect 5181 18173 5215 18207
rect 5549 18173 5583 18207
rect 12909 18173 12943 18207
rect 17417 18173 17451 18207
rect 18337 18173 18371 18207
rect 19257 18173 19291 18207
rect 20545 18173 20579 18207
rect 2881 18105 2915 18139
rect 3709 18105 3743 18139
rect 12725 18105 12759 18139
rect 13645 18105 13679 18139
rect 13829 18105 13863 18139
rect 16313 18105 16347 18139
rect 1501 18037 1535 18071
rect 2007 18037 2041 18071
rect 6101 18037 6135 18071
rect 16865 18037 16899 18071
rect 21557 18037 21591 18071
rect 2559 17833 2593 17867
rect 6929 17833 6963 17867
rect 7481 17833 7515 17867
rect 12265 17833 12299 17867
rect 18061 17833 18095 17867
rect 13185 17765 13219 17799
rect 20177 17765 20211 17799
rect 1777 17697 1811 17731
rect 1961 17697 1995 17731
rect 3065 17697 3099 17731
rect 3341 17697 3375 17731
rect 4169 17697 4203 17731
rect 4445 17697 4479 17731
rect 4905 17697 4939 17731
rect 5089 17697 5123 17731
rect 5825 17697 5859 17731
rect 9873 17697 9907 17731
rect 10149 17697 10183 17731
rect 10517 17697 10551 17731
rect 12541 17697 12575 17731
rect 12909 17697 12943 17731
rect 13369 17697 13403 17731
rect 13829 17697 13863 17731
rect 15577 17697 15611 17731
rect 18337 17697 18371 17731
rect 19257 17697 19291 17731
rect 19533 17697 19567 17731
rect 20729 17697 20763 17731
rect 2053 17629 2087 17663
rect 2630 17629 2664 17663
rect 2973 17629 3007 17663
rect 4077 17629 4111 17663
rect 6009 17629 6043 17663
rect 7113 17629 7147 17663
rect 7389 17629 7423 17663
rect 7665 17629 7699 17663
rect 8953 17629 8987 17663
rect 10241 17629 10275 17663
rect 10609 17629 10643 17663
rect 11069 17629 11103 17663
rect 11345 17629 11379 17663
rect 12449 17629 12483 17663
rect 12817 17629 12851 17663
rect 13461 17629 13495 17663
rect 15393 17629 15427 17663
rect 15485 17629 15519 17663
rect 15853 17629 15887 17663
rect 18429 17629 18463 17663
rect 19625 17629 19659 17663
rect 20545 17629 20579 17663
rect 21154 17629 21188 17663
rect 5181 17561 5215 17595
rect 7297 17561 7331 17595
rect 11161 17561 11195 17595
rect 11529 17561 11563 17595
rect 18889 17561 18923 17595
rect 19073 17561 19107 17595
rect 2421 17493 2455 17527
rect 5549 17493 5583 17527
rect 5917 17493 5951 17527
rect 6377 17493 6411 17527
rect 7573 17493 7607 17527
rect 15025 17493 15059 17527
rect 18705 17493 18739 17527
rect 20637 17493 20671 17527
rect 21051 17493 21085 17527
rect 6009 17289 6043 17323
rect 8861 17289 8895 17323
rect 8953 17289 8987 17323
rect 11069 17289 11103 17323
rect 14289 17289 14323 17323
rect 15117 17289 15151 17323
rect 15577 17289 15611 17323
rect 15853 17289 15887 17323
rect 18797 17289 18831 17323
rect 18889 17289 18923 17323
rect 19349 17289 19383 17323
rect 12633 17221 12667 17255
rect 12817 17221 12851 17255
rect 13001 17221 13035 17255
rect 13829 17221 13863 17255
rect 15209 17221 15243 17255
rect 1685 17153 1719 17187
rect 6193 17153 6227 17187
rect 10425 17153 10459 17187
rect 10885 17153 10919 17187
rect 13277 17153 13311 17187
rect 13461 17153 13495 17187
rect 13921 17153 13955 17187
rect 15669 17153 15703 17187
rect 18613 17153 18647 17187
rect 19073 17153 19107 17187
rect 19533 17153 19567 17187
rect 21373 17153 21407 17187
rect 9045 17085 9079 17119
rect 10057 17085 10091 17119
rect 10517 17085 10551 17119
rect 13093 17085 13127 17119
rect 13645 17085 13679 17119
rect 14933 17085 14967 17119
rect 18429 17085 18463 17119
rect 19717 17085 19751 17119
rect 1501 17017 1535 17051
rect 10701 17017 10735 17051
rect 19257 17017 19291 17051
rect 21557 17017 21591 17051
rect 8493 16949 8527 16983
rect 13001 16745 13035 16779
rect 15669 16745 15703 16779
rect 11161 16677 11195 16711
rect 13093 16677 13127 16711
rect 15577 16677 15611 16711
rect 16497 16677 16531 16711
rect 8309 16609 8343 16643
rect 8401 16609 8435 16643
rect 9965 16609 9999 16643
rect 10517 16609 10551 16643
rect 10701 16609 10735 16643
rect 12449 16609 12483 16643
rect 13645 16609 13679 16643
rect 15761 16609 15795 16643
rect 1409 16541 1443 16575
rect 5641 16541 5675 16575
rect 7205 16541 7239 16575
rect 7757 16541 7791 16575
rect 9660 16541 9694 16575
rect 13461 16541 13495 16575
rect 15853 16541 15887 16575
rect 16313 16541 16347 16575
rect 22017 16541 22051 16575
rect 10793 16473 10827 16507
rect 10977 16473 11011 16507
rect 12633 16473 12667 16507
rect 15393 16473 15427 16507
rect 1593 16405 1627 16439
rect 7021 16405 7055 16439
rect 7573 16405 7607 16439
rect 7849 16405 7883 16439
rect 8217 16405 8251 16439
rect 9505 16405 9539 16439
rect 9873 16405 9907 16439
rect 10333 16405 10367 16439
rect 12541 16405 12575 16439
rect 13553 16405 13587 16439
rect 15485 16405 15519 16439
rect 16037 16405 16071 16439
rect 21833 16405 21867 16439
rect 3985 16201 4019 16235
rect 5733 16201 5767 16235
rect 6837 16201 6871 16235
rect 10609 16201 10643 16235
rect 13047 16201 13081 16235
rect 13415 16201 13449 16235
rect 15301 16201 15335 16235
rect 17233 16201 17267 16235
rect 17693 16201 17727 16235
rect 18061 16201 18095 16235
rect 6745 16133 6779 16167
rect 10977 16133 11011 16167
rect 1685 16065 1719 16099
rect 2421 16065 2455 16099
rect 2605 16065 2639 16099
rect 3341 16065 3375 16099
rect 3617 16065 3651 16099
rect 3801 16065 3835 16099
rect 5641 16065 5675 16099
rect 7021 16065 7055 16099
rect 8677 16065 8711 16099
rect 10400 16065 10434 16099
rect 11069 16065 11103 16099
rect 11575 16065 11609 16099
rect 11678 16065 11712 16099
rect 13150 16065 13184 16099
rect 13486 16065 13520 16099
rect 15669 16065 15703 16099
rect 17601 16065 17635 16099
rect 18429 16065 18463 16099
rect 18521 16065 18555 16099
rect 18889 16065 18923 16099
rect 22017 16065 22051 16099
rect 3157 15997 3191 16031
rect 5825 15997 5859 16031
rect 6377 15997 6411 16031
rect 11253 15997 11287 16031
rect 15761 15997 15795 16031
rect 15853 15997 15887 16031
rect 17785 15997 17819 16031
rect 18613 15997 18647 16031
rect 6561 15929 6595 15963
rect 8861 15929 8895 15963
rect 1501 15861 1535 15895
rect 2789 15861 2823 15895
rect 5273 15861 5307 15895
rect 6469 15861 6503 15895
rect 6745 15861 6779 15895
rect 10471 15861 10505 15895
rect 16221 15861 16255 15895
rect 21833 15861 21867 15895
rect 2421 15657 2455 15691
rect 3249 15657 3283 15691
rect 5917 15657 5951 15691
rect 6285 15657 6319 15691
rect 7757 15657 7791 15691
rect 10517 15657 10551 15691
rect 12449 15657 12483 15691
rect 15761 15657 15795 15691
rect 18429 15657 18463 15691
rect 19533 15657 19567 15691
rect 1869 15521 1903 15555
rect 2697 15521 2731 15555
rect 3893 15521 3927 15555
rect 4077 15521 4111 15555
rect 5365 15521 5399 15555
rect 5457 15521 5491 15555
rect 8401 15521 8435 15555
rect 10977 15521 11011 15555
rect 11069 15521 11103 15555
rect 16221 15521 16255 15555
rect 16313 15521 16347 15555
rect 18889 15521 18923 15555
rect 1409 15453 1443 15487
rect 2881 15453 2915 15487
rect 3474 15453 3508 15487
rect 6469 15453 6503 15487
rect 8585 15453 8619 15487
rect 10885 15453 10919 15487
rect 12633 15453 12667 15487
rect 18797 15453 18831 15487
rect 19257 15453 19291 15487
rect 19349 15453 19383 15487
rect 20520 15453 20554 15487
rect 22017 15453 22051 15487
rect 2053 15385 2087 15419
rect 2789 15385 2823 15419
rect 3387 15385 3421 15419
rect 5549 15385 5583 15419
rect 8217 15385 8251 15419
rect 1593 15317 1627 15351
rect 1961 15317 1995 15351
rect 4169 15317 4203 15351
rect 4537 15317 4571 15351
rect 8125 15317 8159 15351
rect 16129 15317 16163 15351
rect 20591 15317 20625 15351
rect 21833 15317 21867 15351
rect 2099 15113 2133 15147
rect 2881 15113 2915 15147
rect 3985 15113 4019 15147
rect 7757 15113 7791 15147
rect 8217 15113 8251 15147
rect 13001 15113 13035 15147
rect 18337 15113 18371 15147
rect 19901 15113 19935 15147
rect 21097 15113 21131 15147
rect 21189 15113 21223 15147
rect 4445 15045 4479 15079
rect 17877 15045 17911 15079
rect 18245 15045 18279 15079
rect 20269 15045 20303 15079
rect 2028 14977 2062 15011
rect 2697 14977 2731 15011
rect 3157 14977 3191 15011
rect 4905 14977 4939 15011
rect 5273 14977 5307 15011
rect 7481 14977 7515 15011
rect 8125 14977 8159 15011
rect 8953 14977 8987 15011
rect 12633 14977 12667 15011
rect 15945 14977 15979 15011
rect 18061 14977 18095 15011
rect 18705 14977 18739 15011
rect 19533 14977 19567 15011
rect 2513 14909 2547 14943
rect 3065 14909 3099 14943
rect 3525 14909 3559 14943
rect 3801 14909 3835 14943
rect 4997 14909 5031 14943
rect 5181 14909 5215 14943
rect 5641 14909 5675 14943
rect 8309 14909 8343 14943
rect 9045 14909 9079 14943
rect 9137 14909 9171 14943
rect 12449 14909 12483 14943
rect 12541 14909 12575 14943
rect 15853 14909 15887 14943
rect 16313 14909 16347 14943
rect 18797 14909 18831 14943
rect 18889 14909 18923 14943
rect 19165 14909 19199 14943
rect 19625 14909 19659 14943
rect 20361 14909 20395 14943
rect 20453 14909 20487 14943
rect 21281 14909 21315 14943
rect 3617 14841 3651 14875
rect 8585 14841 8619 14875
rect 20729 14841 20763 14875
rect 7665 14773 7699 14807
rect 13461 14773 13495 14807
rect 6101 14569 6135 14603
rect 8953 14569 8987 14603
rect 9413 14569 9447 14603
rect 10149 14569 10183 14603
rect 13093 14569 13127 14603
rect 15485 14569 15519 14603
rect 15577 14569 15611 14603
rect 16497 14569 16531 14603
rect 19257 14569 19291 14603
rect 20407 14569 20441 14603
rect 9781 14501 9815 14535
rect 17877 14501 17911 14535
rect 19625 14501 19659 14535
rect 5549 14433 5583 14467
rect 6745 14433 6779 14467
rect 13553 14433 13587 14467
rect 13737 14433 13771 14467
rect 15209 14433 15243 14467
rect 16129 14433 16163 14467
rect 17509 14433 17543 14467
rect 1409 14365 1443 14399
rect 6653 14365 6687 14399
rect 7021 14365 7055 14399
rect 9137 14365 9171 14399
rect 9597 14365 9631 14399
rect 9873 14365 9907 14399
rect 9965 14365 9999 14399
rect 13001 14365 13035 14399
rect 14657 14365 14691 14399
rect 15117 14365 15151 14399
rect 15945 14365 15979 14399
rect 16957 14365 16991 14399
rect 17417 14365 17451 14399
rect 17693 14365 17727 14399
rect 18705 14365 18739 14399
rect 19441 14365 19475 14399
rect 20510 14365 20544 14399
rect 22017 14365 22051 14399
rect 5641 14297 5675 14331
rect 9321 14297 9355 14331
rect 12633 14297 12667 14331
rect 16037 14297 16071 14331
rect 17049 14297 17083 14331
rect 17233 14297 17267 14331
rect 18889 14297 18923 14331
rect 1593 14229 1627 14263
rect 5733 14229 5767 14263
rect 6193 14229 6227 14263
rect 6561 14229 6595 14263
rect 13461 14229 13495 14263
rect 14197 14229 14231 14263
rect 18521 14229 18555 14263
rect 21833 14229 21867 14263
rect 9873 14025 9907 14059
rect 10241 14025 10275 14059
rect 13001 14025 13035 14059
rect 16497 14025 16531 14059
rect 16681 14025 16715 14059
rect 18613 14025 18647 14059
rect 4629 13957 4663 13991
rect 5457 13957 5491 13991
rect 11989 13957 12023 13991
rect 15669 13957 15703 13991
rect 16313 13957 16347 13991
rect 17049 13957 17083 13991
rect 1409 13889 1443 13923
rect 4445 13889 4479 13923
rect 4813 13889 4847 13923
rect 4997 13889 5031 13923
rect 5365 13889 5399 13923
rect 5917 13889 5951 13923
rect 6009 13889 6043 13923
rect 6745 13889 6779 13923
rect 8677 13889 8711 13923
rect 9137 13889 9171 13923
rect 10333 13889 10367 13923
rect 10747 13889 10781 13923
rect 10850 13889 10884 13923
rect 11094 13889 11128 13923
rect 11805 13889 11839 13923
rect 12173 13889 12207 13923
rect 12541 13889 12575 13923
rect 12633 13889 12667 13923
rect 13737 13889 13771 13923
rect 15393 13889 15427 13923
rect 15577 13889 15611 13923
rect 16129 13889 16163 13923
rect 17141 13889 17175 13923
rect 17555 13889 17589 13923
rect 17658 13889 17692 13923
rect 18797 13889 18831 13923
rect 22017 13889 22051 13923
rect 6377 13821 6411 13855
rect 6653 13821 6687 13855
rect 8309 13821 8343 13855
rect 8769 13821 8803 13855
rect 9229 13821 9263 13855
rect 9505 13821 9539 13855
rect 10517 13821 10551 13855
rect 12449 13821 12483 13855
rect 13369 13821 13403 13855
rect 13645 13821 13679 13855
rect 15209 13821 15243 13855
rect 15853 13821 15887 13855
rect 16037 13821 16071 13855
rect 17233 13821 17267 13855
rect 18981 13821 19015 13855
rect 1593 13753 1627 13787
rect 11023 13685 11057 13719
rect 21833 13685 21867 13719
rect 5457 13481 5491 13515
rect 9781 13481 9815 13515
rect 11345 13481 11379 13515
rect 15301 13481 15335 13515
rect 4629 13413 4663 13447
rect 8953 13413 8987 13447
rect 9873 13413 9907 13447
rect 4353 13345 4387 13379
rect 4813 13345 4847 13379
rect 6009 13345 6043 13379
rect 9137 13345 9171 13379
rect 10333 13345 10367 13379
rect 10517 13345 10551 13379
rect 11529 13345 11563 13379
rect 11713 13345 11747 13379
rect 11989 13345 12023 13379
rect 12725 13345 12759 13379
rect 13185 13345 13219 13379
rect 13921 13345 13955 13379
rect 15853 13345 15887 13379
rect 1409 13277 1443 13311
rect 4261 13277 4295 13311
rect 4997 13277 5031 13311
rect 5549 13277 5583 13311
rect 5733 13277 5767 13311
rect 6193 13277 6227 13311
rect 9597 13277 9631 13311
rect 12817 13277 12851 13311
rect 13829 13277 13863 13311
rect 15669 13277 15703 13311
rect 16246 13277 16280 13311
rect 22017 13277 22051 13311
rect 5089 13209 5123 13243
rect 5917 13209 5951 13243
rect 9321 13209 9355 13243
rect 9413 13209 9447 13243
rect 10241 13209 10275 13243
rect 13369 13209 13403 13243
rect 1593 13141 1627 13175
rect 6377 13141 6411 13175
rect 12081 13141 12115 13175
rect 12173 13141 12207 13175
rect 12541 13141 12575 13175
rect 15761 13141 15795 13175
rect 16175 13141 16209 13175
rect 21833 13141 21867 13175
rect 1593 12937 1627 12971
rect 3893 12937 3927 12971
rect 4261 12937 4295 12971
rect 5181 12937 5215 12971
rect 12127 12937 12161 12971
rect 13001 12937 13035 12971
rect 4721 12869 4755 12903
rect 13829 12869 13863 12903
rect 19625 12869 19659 12903
rect 20453 12869 20487 12903
rect 1409 12801 1443 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 7803 12801 7837 12835
rect 7906 12801 7940 12835
rect 12056 12801 12090 12835
rect 12633 12801 12667 12835
rect 13277 12801 13311 12835
rect 13461 12801 13495 12835
rect 13645 12801 13679 12835
rect 22017 12801 22051 12835
rect 3617 12733 3651 12767
rect 3801 12733 3835 12767
rect 4445 12733 4479 12767
rect 4629 12733 4663 12767
rect 5365 12733 5399 12767
rect 5549 12733 5583 12767
rect 7573 12733 7607 12767
rect 12449 12733 12483 12767
rect 12541 12733 12575 12767
rect 13093 12733 13127 12767
rect 18245 12733 18279 12767
rect 18705 12733 18739 12767
rect 19717 12733 19751 12767
rect 19901 12733 19935 12767
rect 20545 12733 20579 12767
rect 20729 12733 20763 12767
rect 5089 12665 5123 12699
rect 18061 12665 18095 12699
rect 18889 12665 18923 12699
rect 19257 12665 19291 12699
rect 20085 12665 20119 12699
rect 21833 12665 21867 12699
rect 6929 12597 6963 12631
rect 14013 12597 14047 12631
rect 18429 12597 18463 12631
rect 18521 12597 18555 12631
rect 4307 12393 4341 12427
rect 4767 12393 4801 12427
rect 9413 12393 9447 12427
rect 12587 12393 12621 12427
rect 19579 12393 19613 12427
rect 19855 12393 19889 12427
rect 6561 12325 6595 12359
rect 7665 12257 7699 12291
rect 10333 12257 10367 12291
rect 17417 12257 17451 12291
rect 17877 12257 17911 12291
rect 18705 12257 18739 12291
rect 4378 12189 4412 12223
rect 4696 12189 4730 12223
rect 6745 12189 6779 12223
rect 7966 12189 8000 12223
rect 10149 12189 10183 12223
rect 12658 12189 12692 12223
rect 16865 12189 16899 12223
rect 17049 12189 17083 12223
rect 17785 12189 17819 12223
rect 18429 12189 18463 12223
rect 19476 12189 19510 12223
rect 19784 12189 19818 12223
rect 9597 12121 9631 12155
rect 9781 12121 9815 12155
rect 9965 12121 9999 12155
rect 6929 12053 6963 12087
rect 7021 12053 7055 12087
rect 7389 12053 7423 12087
rect 7481 12053 7515 12087
rect 7895 12053 7929 12087
rect 17141 12053 17175 12087
rect 18061 12053 18095 12087
rect 18521 12053 18555 12087
rect 7113 11849 7147 11883
rect 8953 11849 8987 11883
rect 17141 11849 17175 11883
rect 17509 11849 17543 11883
rect 17969 11849 18003 11883
rect 18337 11849 18371 11883
rect 7205 11781 7239 11815
rect 8401 11781 8435 11815
rect 15761 11781 15795 11815
rect 16037 11781 16071 11815
rect 17049 11781 17083 11815
rect 18521 11781 18555 11815
rect 18705 11781 18739 11815
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 2088 11713 2122 11747
rect 7757 11713 7791 11747
rect 8033 11713 8067 11747
rect 8217 11713 8251 11747
rect 9229 11713 9263 11747
rect 10241 11713 10275 11747
rect 11529 11713 11563 11747
rect 14289 11713 14323 11747
rect 15301 11713 15335 11747
rect 15853 11713 15887 11747
rect 17877 11713 17911 11747
rect 22017 11713 22051 11747
rect 7297 11645 7331 11679
rect 8769 11645 8803 11679
rect 9137 11645 9171 11679
rect 9873 11645 9907 11679
rect 10333 11645 10367 11679
rect 10701 11645 10735 11679
rect 14197 11645 14231 11679
rect 15393 11645 15427 11679
rect 15577 11645 15611 11679
rect 17233 11645 17267 11679
rect 18061 11645 18095 11679
rect 1593 11577 1627 11611
rect 1869 11577 1903 11611
rect 7941 11577 7975 11611
rect 8585 11577 8619 11611
rect 10885 11577 10919 11611
rect 21833 11577 21867 11611
rect 2191 11509 2225 11543
rect 6745 11509 6779 11543
rect 7573 11509 7607 11543
rect 9597 11509 9631 11543
rect 10517 11509 10551 11543
rect 11713 11509 11747 11543
rect 14657 11509 14691 11543
rect 14841 11509 14875 11543
rect 16221 11509 16255 11543
rect 16681 11509 16715 11543
rect 8033 11305 8067 11339
rect 11989 11305 12023 11339
rect 13921 11305 13955 11339
rect 18153 11305 18187 11339
rect 11161 11237 11195 11271
rect 17417 11237 17451 11271
rect 18245 11237 18279 11271
rect 21833 11237 21867 11271
rect 6929 11169 6963 11203
rect 7205 11169 7239 11203
rect 9689 11169 9723 11203
rect 10793 11169 10827 11203
rect 11805 11169 11839 11203
rect 12541 11169 12575 11203
rect 13553 11169 13587 11203
rect 13737 11169 13771 11203
rect 14197 11169 14231 11203
rect 15577 11169 15611 11203
rect 16957 11169 16991 11203
rect 17693 11169 17727 11203
rect 18429 11169 18463 11203
rect 1501 11101 1535 11135
rect 2697 11101 2731 11135
rect 2881 11101 2915 11135
rect 3525 11101 3559 11135
rect 5089 11101 5123 11135
rect 6837 11101 6871 11135
rect 7665 11101 7699 11135
rect 9413 11101 9447 11135
rect 9505 11101 9539 11135
rect 9873 11101 9907 11135
rect 10609 11101 10643 11135
rect 13328 11101 13362 11135
rect 14381 11101 14415 11135
rect 14473 11101 14507 11135
rect 15910 11101 15944 11135
rect 17785 11101 17819 11135
rect 18613 11101 18647 11135
rect 18889 11101 18923 11135
rect 22017 11101 22051 11135
rect 1961 11033 1995 11067
rect 3065 11033 3099 11067
rect 4537 11033 4571 11067
rect 4721 11033 4755 11067
rect 4905 11033 4939 11067
rect 7849 11033 7883 11067
rect 12449 11033 12483 11067
rect 13415 11033 13449 11067
rect 15301 11033 15335 11067
rect 15393 11033 15427 11067
rect 15807 11033 15841 11067
rect 18705 11033 18739 11067
rect 1685 10965 1719 10999
rect 3249 10965 3283 10999
rect 3433 10965 3467 10999
rect 9045 10965 9079 10999
rect 10241 10965 10275 10999
rect 10701 10965 10735 10999
rect 11529 10965 11563 10999
rect 11621 10965 11655 10999
rect 12357 10965 12391 10999
rect 14841 10965 14875 10999
rect 14933 10965 14967 10999
rect 19073 10965 19107 10999
rect 1593 10761 1627 10795
rect 3157 10761 3191 10795
rect 5181 10761 5215 10795
rect 9229 10761 9263 10795
rect 11667 10761 11701 10795
rect 12035 10761 12069 10795
rect 2421 10693 2455 10727
rect 5917 10693 5951 10727
rect 7941 10693 7975 10727
rect 9137 10693 9171 10727
rect 11345 10693 11379 10727
rect 15117 10693 15151 10727
rect 1777 10625 1811 10659
rect 3249 10625 3283 10659
rect 3893 10625 3927 10659
rect 5089 10625 5123 10659
rect 6929 10625 6963 10659
rect 7481 10625 7515 10659
rect 11738 10625 11772 10659
rect 11932 10625 11966 10659
rect 14473 10625 14507 10659
rect 14933 10625 14967 10659
rect 19257 10625 19291 10659
rect 19441 10625 19475 10659
rect 19901 10625 19935 10659
rect 20510 10625 20544 10659
rect 22017 10625 22051 10659
rect 2237 10557 2271 10591
rect 2329 10557 2363 10591
rect 2973 10557 3007 10591
rect 3801 10557 3835 10591
rect 5365 10557 5399 10591
rect 7021 10557 7055 10591
rect 7389 10557 7423 10591
rect 9413 10557 9447 10591
rect 14013 10557 14047 10591
rect 14565 10557 14599 10591
rect 19717 10557 19751 10591
rect 1961 10489 1995 10523
rect 2789 10489 2823 10523
rect 3617 10489 3651 10523
rect 13829 10489 13863 10523
rect 14841 10489 14875 10523
rect 21833 10489 21867 10523
rect 4261 10421 4295 10455
rect 4721 10421 4755 10455
rect 5825 10421 5859 10455
rect 7297 10421 7331 10455
rect 8769 10421 8803 10455
rect 10057 10421 10091 10455
rect 14197 10421 14231 10455
rect 15301 10421 15335 10455
rect 19625 10421 19659 10455
rect 20085 10421 20119 10455
rect 20407 10421 20441 10455
rect 2835 10217 2869 10251
rect 3433 10217 3467 10251
rect 4537 10217 4571 10251
rect 8309 10217 8343 10251
rect 10793 10217 10827 10251
rect 12265 10217 12299 10251
rect 20085 10217 20119 10251
rect 2697 10149 2731 10183
rect 3065 10149 3099 10183
rect 5365 10149 5399 10183
rect 12449 10149 12483 10183
rect 16681 10149 16715 10183
rect 2145 10081 2179 10115
rect 2237 10081 2271 10115
rect 3249 10081 3283 10115
rect 4261 10081 4295 10115
rect 4813 10081 4847 10115
rect 4905 10081 4939 10115
rect 14473 10081 14507 10115
rect 14565 10081 14599 10115
rect 17417 10081 17451 10115
rect 18337 10081 18371 10115
rect 18521 10081 18555 10115
rect 19717 10081 19751 10115
rect 19809 10081 19843 10115
rect 20545 10081 20579 10115
rect 20637 10081 20671 10115
rect 21465 10081 21499 10115
rect 1685 10013 1719 10047
rect 2329 10013 2363 10047
rect 2906 10013 2940 10047
rect 4169 10013 4203 10047
rect 4997 10013 5031 10047
rect 5641 10013 5675 10047
rect 6653 10013 6687 10047
rect 6929 10013 6963 10047
rect 10425 10013 10459 10047
rect 10609 10013 10643 10047
rect 12081 10013 12115 10047
rect 12265 10013 12299 10047
rect 12357 10013 12391 10047
rect 12560 10013 12594 10047
rect 12725 10013 12759 10047
rect 12817 10013 12851 10047
rect 13185 10013 13219 10047
rect 14657 10013 14691 10047
rect 16497 10013 16531 10047
rect 20453 10013 20487 10047
rect 21741 10013 21775 10047
rect 7021 9945 7055 9979
rect 13093 9945 13127 9979
rect 17233 9945 17267 9979
rect 1501 9877 1535 9911
rect 5457 9877 5491 9911
rect 6469 9877 6503 9911
rect 12449 9877 12483 9911
rect 12817 9877 12851 9911
rect 13001 9877 13035 9911
rect 15025 9877 15059 9911
rect 16865 9877 16899 9911
rect 17325 9877 17359 9911
rect 17693 9877 17727 9911
rect 18061 9877 18095 9911
rect 18153 9877 18187 9911
rect 18981 9877 19015 9911
rect 19257 9877 19291 9911
rect 19625 9877 19659 9911
rect 20913 9877 20947 9911
rect 21281 9877 21315 9911
rect 21373 9877 21407 9911
rect 21925 9877 21959 9911
rect 16773 9673 16807 9707
rect 20637 9673 20671 9707
rect 20867 9673 20901 9707
rect 4813 9605 4847 9639
rect 7849 9605 7883 9639
rect 15209 9605 15243 9639
rect 20177 9605 20211 9639
rect 4353 9537 4387 9571
rect 6653 9537 6687 9571
rect 6837 9537 6871 9571
rect 7205 9537 7239 9571
rect 7757 9537 7791 9571
rect 15025 9537 15059 9571
rect 16313 9537 16347 9571
rect 16773 9537 16807 9571
rect 17141 9537 17175 9571
rect 17417 9537 17451 9571
rect 17877 9537 17911 9571
rect 18245 9537 18279 9571
rect 18889 9537 18923 9571
rect 19533 9537 19567 9571
rect 19993 9537 20027 9571
rect 20796 9537 20830 9571
rect 4261 9469 4295 9503
rect 18521 9469 18555 9503
rect 18797 9469 18831 9503
rect 19165 9469 19199 9503
rect 19441 9469 19475 9503
rect 20269 9469 20303 9503
rect 20453 9469 20487 9503
rect 16497 9401 16531 9435
rect 15485 9333 15519 9367
rect 19809 9333 19843 9367
rect 6745 9129 6779 9163
rect 18797 9129 18831 9163
rect 1501 9061 1535 9095
rect 7665 9061 7699 9095
rect 15025 9061 15059 9095
rect 18429 9061 18463 9095
rect 6193 8993 6227 9027
rect 7389 8993 7423 9027
rect 14381 8993 14415 9027
rect 15577 8993 15611 9027
rect 15669 8993 15703 9027
rect 18613 8993 18647 9027
rect 1685 8925 1719 8959
rect 6377 8925 6411 8959
rect 7205 8925 7239 8959
rect 7849 8925 7883 8959
rect 8953 8925 8987 8959
rect 9413 8925 9447 8959
rect 9597 8925 9631 8959
rect 9689 8925 9723 8959
rect 10368 8925 10402 8959
rect 11069 8925 11103 8959
rect 11253 8925 11287 8959
rect 11345 8925 11379 8959
rect 11846 8925 11880 8959
rect 12541 8925 12575 8959
rect 12633 8925 12667 8959
rect 12817 8925 12851 8959
rect 13369 8925 13403 8959
rect 14657 8925 14691 8959
rect 15485 8925 15519 8959
rect 15945 8925 15979 8959
rect 21741 8925 21775 8959
rect 6285 8857 6319 8891
rect 10609 8857 10643 8891
rect 11759 8857 11793 8891
rect 13277 8857 13311 8891
rect 14565 8857 14599 8891
rect 6837 8789 6871 8823
rect 7297 8789 7331 8823
rect 10471 8789 10505 8823
rect 15117 8789 15151 8823
rect 16129 8789 16163 8823
rect 21925 8789 21959 8823
rect 4445 8585 4479 8619
rect 8401 8585 8435 8619
rect 9229 8585 9263 8619
rect 9597 8585 9631 8619
rect 3157 8517 3191 8551
rect 11529 8517 11563 8551
rect 12725 8517 12759 8551
rect 1685 8449 1719 8483
rect 2789 8449 2823 8483
rect 2973 8449 3007 8483
rect 3433 8449 3467 8483
rect 4077 8449 4111 8483
rect 4261 8449 4295 8483
rect 4813 8449 4847 8483
rect 8217 8449 8251 8483
rect 9781 8449 9815 8483
rect 11989 8449 12023 8483
rect 12173 8449 12207 8483
rect 13185 8449 13219 8483
rect 13369 8449 13403 8483
rect 14657 8449 14691 8483
rect 16681 8449 16715 8483
rect 19993 8449 20027 8483
rect 21373 8449 21407 8483
rect 4721 8381 4755 8415
rect 8585 8381 8619 8415
rect 9045 8381 9079 8415
rect 9137 8381 9171 8415
rect 10793 8381 10827 8415
rect 12265 8381 12299 8415
rect 13461 8381 13495 8415
rect 19165 8381 19199 8415
rect 19349 8381 19383 8415
rect 1501 8313 1535 8347
rect 3249 8313 3283 8347
rect 3617 8313 3651 8347
rect 5181 8313 5215 8347
rect 8033 8313 8067 8347
rect 8769 8313 8803 8347
rect 14841 8313 14875 8347
rect 16865 8313 16899 8347
rect 21557 8313 21591 8347
rect 5641 8245 5675 8279
rect 17601 8245 17635 8279
rect 18981 8245 19015 8279
rect 19533 8245 19567 8279
rect 3065 8041 3099 8075
rect 3525 8041 3559 8075
rect 9137 8041 9171 8075
rect 11713 8041 11747 8075
rect 12633 8041 12667 8075
rect 2237 7973 2271 8007
rect 8217 7973 8251 8007
rect 15853 7973 15887 8007
rect 1685 7905 1719 7939
rect 2513 7905 2547 7939
rect 3157 7905 3191 7939
rect 3341 7905 3375 7939
rect 3985 7905 4019 7939
rect 4077 7905 4111 7939
rect 5641 7905 5675 7939
rect 5733 7905 5767 7939
rect 8033 7905 8067 7939
rect 9597 7905 9631 7939
rect 11069 7905 11103 7939
rect 11253 7905 11287 7939
rect 11805 7905 11839 7939
rect 13277 7905 13311 7939
rect 14565 7905 14599 7939
rect 16957 7905 16991 7939
rect 17693 7905 17727 7939
rect 17785 7905 17819 7939
rect 18521 7905 18555 7939
rect 18981 7905 19015 7939
rect 19809 7905 19843 7939
rect 4169 7837 4203 7871
rect 5549 7837 5583 7871
rect 6653 7837 6687 7871
rect 7205 7837 7239 7871
rect 7941 7837 7975 7871
rect 8217 7837 8251 7871
rect 9321 7837 9355 7871
rect 9505 7837 9539 7871
rect 9781 7837 9815 7871
rect 10333 7837 10367 7871
rect 10425 7837 10459 7871
rect 10609 7837 10643 7871
rect 11345 7837 11379 7871
rect 11989 7837 12023 7871
rect 14749 7837 14783 7871
rect 14841 7837 14875 7871
rect 15117 7837 15151 7871
rect 15301 7837 15335 7871
rect 15669 7837 15703 7871
rect 18889 7837 18923 7871
rect 21741 7837 21775 7871
rect 7849 7769 7883 7803
rect 16773 7769 16807 7803
rect 17601 7769 17635 7803
rect 1777 7701 1811 7735
rect 1869 7701 1903 7735
rect 2605 7701 2639 7735
rect 2697 7701 2731 7735
rect 4537 7701 4571 7735
rect 5181 7701 5215 7735
rect 6469 7701 6503 7735
rect 7389 7701 7423 7735
rect 9965 7701 9999 7735
rect 12173 7701 12207 7735
rect 13001 7701 13035 7735
rect 13093 7701 13127 7735
rect 16405 7701 16439 7735
rect 16865 7701 16899 7735
rect 17233 7701 17267 7735
rect 19257 7701 19291 7735
rect 19625 7701 19659 7735
rect 19717 7701 19751 7735
rect 21925 7701 21959 7735
rect 1593 7497 1627 7531
rect 2099 7497 2133 7531
rect 2743 7497 2777 7531
rect 5365 7497 5399 7531
rect 5825 7497 5859 7531
rect 13185 7497 13219 7531
rect 18797 7497 18831 7531
rect 4445 7429 4479 7463
rect 5457 7429 5491 7463
rect 9965 7429 9999 7463
rect 10149 7429 10183 7463
rect 12725 7429 12759 7463
rect 18521 7429 18555 7463
rect 20637 7429 20671 7463
rect 1409 7361 1443 7395
rect 1685 7361 1719 7395
rect 2170 7361 2204 7395
rect 2640 7361 2674 7395
rect 3249 7361 3283 7395
rect 4905 7361 4939 7395
rect 7665 7361 7699 7395
rect 12375 7361 12409 7395
rect 12541 7361 12575 7395
rect 13001 7361 13035 7395
rect 14473 7361 14507 7395
rect 15117 7361 15151 7395
rect 18705 7361 18739 7395
rect 19625 7361 19659 7395
rect 20729 7361 20763 7395
rect 21143 7361 21177 7395
rect 21246 7361 21280 7395
rect 21522 7361 21556 7395
rect 22017 7361 22051 7395
rect 3157 7293 3191 7327
rect 3617 7293 3651 7327
rect 4997 7293 5031 7327
rect 5273 7293 5307 7327
rect 12817 7293 12851 7327
rect 18981 7293 19015 7327
rect 19165 7293 19199 7327
rect 19257 7293 19291 7327
rect 19533 7293 19567 7327
rect 20821 7293 20855 7327
rect 1869 7225 1903 7259
rect 14657 7225 14691 7259
rect 20269 7225 20303 7259
rect 21833 7225 21867 7259
rect 7849 7157 7883 7191
rect 10333 7157 10367 7191
rect 15301 7157 15335 7191
rect 18337 7157 18371 7191
rect 21419 7157 21453 7191
rect 6561 6953 6595 6987
rect 15577 6953 15611 6987
rect 19901 6953 19935 6987
rect 20453 6885 20487 6919
rect 6009 6817 6043 6851
rect 12633 6817 12667 6851
rect 13093 6817 13127 6851
rect 16129 6817 16163 6851
rect 17417 6817 17451 6851
rect 18245 6817 18279 6851
rect 19257 6817 19291 6851
rect 20913 6817 20947 6851
rect 21005 6817 21039 6851
rect 5457 6749 5491 6783
rect 6837 6749 6871 6783
rect 8401 6749 8435 6783
rect 13001 6749 13035 6783
rect 18153 6749 18187 6783
rect 18521 6749 18555 6783
rect 20085 6749 20119 6783
rect 20269 6749 20303 6783
rect 5089 6681 5123 6715
rect 6193 6681 6227 6715
rect 15945 6681 15979 6715
rect 17233 6681 17267 6715
rect 6101 6613 6135 6647
rect 8585 6613 8619 6647
rect 16037 6613 16071 6647
rect 16865 6613 16899 6647
rect 17325 6613 17359 6647
rect 17693 6613 17727 6647
rect 18061 6613 18095 6647
rect 19717 6613 19751 6647
rect 20821 6613 20855 6647
rect 1593 6409 1627 6443
rect 4445 6409 4479 6443
rect 5273 6409 5307 6443
rect 6377 6409 6411 6443
rect 6837 6409 6871 6443
rect 8033 6409 8067 6443
rect 8861 6409 8895 6443
rect 9321 6409 9355 6443
rect 9689 6409 9723 6443
rect 16681 6409 16715 6443
rect 19901 6409 19935 6443
rect 4261 6341 4295 6375
rect 5457 6341 5491 6375
rect 14657 6341 14691 6375
rect 14749 6341 14783 6375
rect 1409 6273 1443 6307
rect 3744 6273 3778 6307
rect 4077 6273 4111 6307
rect 4905 6273 4939 6307
rect 6745 6273 6779 6307
rect 7665 6273 7699 6307
rect 9229 6273 9263 6307
rect 10057 6273 10091 6307
rect 10149 6273 10183 6307
rect 10517 6273 10551 6307
rect 12357 6273 12391 6307
rect 13001 6273 13035 6307
rect 13461 6273 13495 6307
rect 17049 6273 17083 6307
rect 18797 6273 18831 6307
rect 20085 6273 20119 6307
rect 21373 6273 21407 6307
rect 4721 6205 4755 6239
rect 4813 6205 4847 6239
rect 5733 6205 5767 6239
rect 7021 6205 7055 6239
rect 7481 6205 7515 6239
rect 7573 6205 7607 6239
rect 9413 6205 9447 6239
rect 10241 6205 10275 6239
rect 11897 6205 11931 6239
rect 12449 6205 12483 6239
rect 12725 6205 12759 6239
rect 12817 6205 12851 6239
rect 13553 6205 13587 6239
rect 14565 6205 14599 6239
rect 16497 6205 16531 6239
rect 17141 6205 17175 6239
rect 17233 6205 17267 6239
rect 18429 6205 18463 6239
rect 18889 6205 18923 6239
rect 20269 6205 20303 6239
rect 12081 6137 12115 6171
rect 14197 6137 14231 6171
rect 21557 6137 21591 6171
rect 3847 6069 3881 6103
rect 8125 6069 8159 6103
rect 11713 6069 11747 6103
rect 13185 6069 13219 6103
rect 13829 6069 13863 6103
rect 14933 6069 14967 6103
rect 3249 5865 3283 5899
rect 6101 5865 6135 5899
rect 7573 5865 7607 5899
rect 9781 5865 9815 5899
rect 10701 5865 10735 5899
rect 11897 5865 11931 5899
rect 14473 5865 14507 5899
rect 21833 5865 21867 5899
rect 3617 5797 3651 5831
rect 4537 5797 4571 5831
rect 19073 5797 19107 5831
rect 3893 5729 3927 5763
rect 4905 5729 4939 5763
rect 5181 5729 5215 5763
rect 5641 5729 5675 5763
rect 8033 5729 8067 5763
rect 8217 5729 8251 5763
rect 10057 5729 10091 5763
rect 10425 5729 10459 5763
rect 12449 5729 12483 5763
rect 14933 5729 14967 5763
rect 15025 5729 15059 5763
rect 1685 5661 1719 5695
rect 3433 5661 3467 5695
rect 4077 5661 4111 5695
rect 4813 5661 4847 5695
rect 5733 5661 5767 5695
rect 10149 5661 10183 5695
rect 10517 5661 10551 5695
rect 11688 5661 11722 5695
rect 12842 5661 12876 5695
rect 13001 5661 13035 5695
rect 13185 5661 13219 5695
rect 18889 5661 18923 5695
rect 22017 5661 22051 5695
rect 12265 5593 12299 5627
rect 1501 5525 1535 5559
rect 4169 5525 4203 5559
rect 7941 5525 7975 5559
rect 11759 5525 11793 5559
rect 12357 5525 12391 5559
rect 12771 5525 12805 5559
rect 13369 5525 13403 5559
rect 14841 5525 14875 5559
rect 18705 5525 18739 5559
rect 1593 5321 1627 5355
rect 4261 5321 4295 5355
rect 4721 5321 4755 5355
rect 11989 5321 12023 5355
rect 12449 5321 12483 5355
rect 18245 5321 18279 5355
rect 21833 5321 21867 5355
rect 4353 5253 4387 5287
rect 4997 5253 5031 5287
rect 7021 5253 7055 5287
rect 8401 5253 8435 5287
rect 9781 5253 9815 5287
rect 1409 5185 1443 5219
rect 4537 5185 4571 5219
rect 5457 5185 5491 5219
rect 6837 5185 6871 5219
rect 7573 5185 7607 5219
rect 9597 5185 9631 5219
rect 12081 5185 12115 5219
rect 14381 5185 14415 5219
rect 16865 5185 16899 5219
rect 18613 5185 18647 5219
rect 19441 5185 19475 5219
rect 22017 5185 22051 5219
rect 3893 5117 3927 5151
rect 4077 5117 4111 5151
rect 5549 5117 5583 5151
rect 7205 5117 7239 5151
rect 7481 5117 7515 5151
rect 7941 5117 7975 5151
rect 8217 5117 8251 5151
rect 9965 5117 9999 5151
rect 11897 5117 11931 5151
rect 13921 5117 13955 5151
rect 14473 5117 14507 5151
rect 16773 5117 16807 5151
rect 17233 5117 17267 5151
rect 17877 5117 17911 5151
rect 18705 5117 18739 5151
rect 18797 5117 18831 5151
rect 19073 5117 19107 5151
rect 19349 5117 19383 5151
rect 8033 5049 8067 5083
rect 17417 5049 17451 5083
rect 1593 4777 1627 4811
rect 9045 4777 9079 4811
rect 10333 4777 10367 4811
rect 13921 4777 13955 4811
rect 15117 4777 15151 4811
rect 17693 4777 17727 4811
rect 18981 4777 19015 4811
rect 19257 4777 19291 4811
rect 9505 4709 9539 4743
rect 17325 4709 17359 4743
rect 18061 4709 18095 4743
rect 18153 4709 18187 4743
rect 5825 4641 5859 4675
rect 7021 4641 7055 4675
rect 9413 4641 9447 4675
rect 10149 4641 10183 4675
rect 10793 4641 10827 4675
rect 14473 4641 14507 4675
rect 15577 4641 15611 4675
rect 16865 4641 16899 4675
rect 18337 4641 18371 4675
rect 20637 4641 20671 4675
rect 1409 4573 1443 4607
rect 5641 4573 5675 4607
rect 7205 4573 7239 4607
rect 9229 4573 9263 4607
rect 10701 4573 10735 4607
rect 13737 4573 13771 4607
rect 15485 4573 15519 4607
rect 15853 4573 15887 4607
rect 16681 4573 16715 4607
rect 17877 4573 17911 4607
rect 18797 4573 18831 4607
rect 19625 4573 19659 4607
rect 20361 4573 20395 4607
rect 20970 4573 21004 4607
rect 22017 4573 22051 4607
rect 9873 4505 9907 4539
rect 13553 4505 13587 4539
rect 16957 4505 16991 4539
rect 17141 4505 17175 4539
rect 18521 4505 18555 4539
rect 18613 4505 18647 4539
rect 19441 4505 19475 4539
rect 7389 4437 7423 4471
rect 9965 4437 9999 4471
rect 14933 4437 14967 4471
rect 15945 4437 15979 4471
rect 16497 4437 16531 4471
rect 19993 4437 20027 4471
rect 20453 4437 20487 4471
rect 20867 4437 20901 4471
rect 21833 4437 21867 4471
rect 4077 4233 4111 4267
rect 7481 4233 7515 4267
rect 10057 4233 10091 4267
rect 10149 4233 10183 4267
rect 13277 4233 13311 4267
rect 14381 4233 14415 4267
rect 18797 4233 18831 4267
rect 4445 4165 4479 4199
rect 5733 4165 5767 4199
rect 19165 4165 19199 4199
rect 4905 4097 4939 4131
rect 6126 4097 6160 4131
rect 6653 4097 6687 4131
rect 9689 4097 9723 4131
rect 9873 4097 9907 4131
rect 11897 4097 11931 4131
rect 13553 4097 13587 4131
rect 15669 4097 15703 4131
rect 15853 4097 15887 4131
rect 16129 4097 16163 4131
rect 17049 4097 17083 4131
rect 4537 4029 4571 4063
rect 4721 4029 4755 4063
rect 6745 4029 6779 4063
rect 7205 4029 7239 4063
rect 7389 4029 7423 4063
rect 10333 4029 10367 4063
rect 11989 4029 12023 4063
rect 12081 4029 12115 4063
rect 12909 4029 12943 4063
rect 13093 4029 13127 4063
rect 13645 4029 13679 4063
rect 14105 4029 14139 4063
rect 14289 4029 14323 4063
rect 16221 4029 16255 4063
rect 16497 4029 16531 4063
rect 17141 4029 17175 4063
rect 17325 4029 17359 4063
rect 19257 4029 19291 4063
rect 19441 4029 19475 4063
rect 6055 3961 6089 3995
rect 7021 3961 7055 3995
rect 7849 3961 7883 3995
rect 10517 3961 10551 3995
rect 11529 3961 11563 3995
rect 14749 3961 14783 3995
rect 15485 3961 15519 3995
rect 13921 3893 13955 3927
rect 16681 3893 16715 3927
rect 1593 3689 1627 3723
rect 5825 3689 5859 3723
rect 7389 3689 7423 3723
rect 9413 3689 9447 3723
rect 11483 3689 11517 3723
rect 13461 3689 13495 3723
rect 13921 3689 13955 3723
rect 16589 3689 16623 3723
rect 17049 3689 17083 3723
rect 19303 3689 19337 3723
rect 6009 3553 6043 3587
rect 6193 3553 6227 3587
rect 10057 3553 10091 3587
rect 13093 3553 13127 3587
rect 16221 3553 16255 3587
rect 16681 3553 16715 3587
rect 7205 3485 7239 3519
rect 11412 3485 11446 3519
rect 13277 3485 13311 3519
rect 14222 3485 14256 3519
rect 16405 3485 16439 3519
rect 16865 3485 16899 3519
rect 17208 3485 17242 3519
rect 19406 3485 19440 3519
rect 1501 3417 1535 3451
rect 7021 3417 7055 3451
rect 9781 3417 9815 3451
rect 13553 3417 13587 3451
rect 13737 3417 13771 3451
rect 14749 3417 14783 3451
rect 9873 3349 9907 3383
rect 14151 3349 14185 3383
rect 14473 3349 14507 3383
rect 17279 3349 17313 3383
rect 7113 3145 7147 3179
rect 9827 3145 9861 3179
rect 13829 3145 13863 3179
rect 14289 3145 14323 3179
rect 14657 3145 14691 3179
rect 16681 3145 16715 3179
rect 17509 3145 17543 3179
rect 17969 3145 18003 3179
rect 7481 3077 7515 3111
rect 6904 3009 6938 3043
rect 7573 3009 7607 3043
rect 7987 3009 8021 3043
rect 8090 3009 8124 3043
rect 9930 3009 9964 3043
rect 13620 3009 13654 3043
rect 14197 3009 14231 3043
rect 15025 3009 15059 3043
rect 16364 3009 16398 3043
rect 17049 3009 17083 3043
rect 17877 3009 17911 3043
rect 7757 2941 7791 2975
rect 14473 2941 14507 2975
rect 15117 2941 15151 2975
rect 15301 2941 15335 2975
rect 16451 2941 16485 2975
rect 17141 2941 17175 2975
rect 17233 2941 17267 2975
rect 18153 2941 18187 2975
rect 13691 2873 13725 2907
rect 6975 2805 7009 2839
rect 4813 2601 4847 2635
rect 5457 2601 5491 2635
rect 6561 2601 6595 2635
rect 9965 2601 9999 2635
rect 10425 2601 10459 2635
rect 11253 2601 11287 2635
rect 11713 2601 11747 2635
rect 12541 2601 12575 2635
rect 14933 2601 14967 2635
rect 18153 2601 18187 2635
rect 19441 2601 19475 2635
rect 20085 2601 20119 2635
rect 3525 2533 3559 2567
rect 4169 2533 4203 2567
rect 9321 2533 9355 2567
rect 13645 2533 13679 2567
rect 17509 2533 17543 2567
rect 7113 2465 7147 2499
rect 7297 2465 7331 2499
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 6193 2397 6227 2431
rect 6377 2397 6411 2431
rect 7481 2397 7515 2431
rect 7849 2397 7883 2431
rect 8493 2397 8527 2431
rect 9137 2397 9171 2431
rect 9781 2397 9815 2431
rect 10609 2397 10643 2431
rect 11069 2397 11103 2431
rect 11897 2397 11931 2431
rect 12357 2397 12391 2431
rect 13001 2397 13035 2431
rect 13829 2397 13863 2431
rect 14289 2397 14323 2431
rect 15117 2397 15151 2431
rect 15577 2397 15611 2431
rect 16221 2397 16255 2431
rect 16865 2397 16899 2431
rect 17693 2397 17727 2431
rect 18337 2397 18371 2431
rect 18797 2397 18831 2431
rect 19625 2397 19659 2431
rect 20269 2397 20303 2431
rect 7021 2329 7055 2363
rect 13277 2329 13311 2363
rect 6009 2261 6043 2295
rect 6653 2261 6687 2295
rect 7665 2261 7699 2295
rect 8033 2261 8067 2295
rect 8677 2261 8711 2295
rect 14473 2261 14507 2295
rect 15761 2261 15795 2295
rect 16405 2261 16439 2295
rect 17049 2261 17083 2295
rect 18981 2261 19015 2295
<< metal1 >>
rect 1104 23418 22356 23440
rect 1104 23366 3606 23418
rect 3658 23366 3670 23418
rect 3722 23366 3734 23418
rect 3786 23366 3798 23418
rect 3850 23366 3862 23418
rect 3914 23366 8919 23418
rect 8971 23366 8983 23418
rect 9035 23366 9047 23418
rect 9099 23366 9111 23418
rect 9163 23366 9175 23418
rect 9227 23366 14232 23418
rect 14284 23366 14296 23418
rect 14348 23366 14360 23418
rect 14412 23366 14424 23418
rect 14476 23366 14488 23418
rect 14540 23366 19545 23418
rect 19597 23366 19609 23418
rect 19661 23366 19673 23418
rect 19725 23366 19737 23418
rect 19789 23366 19801 23418
rect 19853 23366 22356 23418
rect 1104 23344 22356 23366
rect 7098 23264 7104 23316
rect 7156 23304 7162 23316
rect 7377 23307 7435 23313
rect 7377 23304 7389 23307
rect 7156 23276 7389 23304
rect 7156 23264 7162 23276
rect 7377 23273 7389 23276
rect 7423 23273 7435 23307
rect 7377 23267 7435 23273
rect 8018 23264 8024 23316
rect 8076 23264 8082 23316
rect 11606 23264 11612 23316
rect 11664 23264 11670 23316
rect 14090 23264 14096 23316
rect 14148 23304 14154 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 14148 23276 14473 23304
rect 14148 23264 14154 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 16758 23264 16764 23316
rect 16816 23304 16822 23316
rect 17405 23307 17463 23313
rect 17405 23304 17417 23307
rect 16816 23276 17417 23304
rect 16816 23264 16822 23276
rect 17405 23273 17417 23276
rect 17451 23273 17463 23307
rect 17405 23267 17463 23273
rect 18322 23264 18328 23316
rect 18380 23264 18386 23316
rect 9309 23239 9367 23245
rect 9309 23205 9321 23239
rect 9355 23236 9367 23239
rect 11054 23236 11060 23248
rect 9355 23208 11060 23236
rect 9355 23205 9367 23208
rect 9309 23199 9367 23205
rect 11054 23196 11060 23208
rect 11112 23196 11118 23248
rect 12250 23196 12256 23248
rect 12308 23196 12314 23248
rect 16114 23196 16120 23248
rect 16172 23236 16178 23248
rect 16945 23239 17003 23245
rect 16945 23236 16957 23239
rect 16172 23208 16957 23236
rect 16172 23196 16178 23208
rect 16945 23205 16957 23208
rect 16991 23205 17003 23239
rect 16945 23199 17003 23205
rect 18785 23239 18843 23245
rect 18785 23205 18797 23239
rect 18831 23205 18843 23239
rect 18785 23199 18843 23205
rect 13173 23171 13231 23177
rect 13173 23168 13185 23171
rect 11164 23140 13185 23168
rect 4798 23060 4804 23112
rect 4856 23060 4862 23112
rect 5258 23060 5264 23112
rect 5316 23060 5322 23112
rect 6546 23060 6552 23112
rect 6604 23060 6610 23112
rect 8386 23060 8392 23112
rect 8444 23100 8450 23112
rect 8665 23103 8723 23109
rect 8665 23100 8677 23103
rect 8444 23072 8677 23100
rect 8444 23060 8450 23072
rect 8665 23069 8677 23072
rect 8711 23069 8723 23103
rect 8665 23063 8723 23069
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9306 23100 9312 23112
rect 9171 23072 9312 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9306 23060 9312 23072
rect 9364 23060 9370 23112
rect 9674 23060 9680 23112
rect 9732 23100 9738 23112
rect 9769 23103 9827 23109
rect 9769 23100 9781 23103
rect 9732 23072 9781 23100
rect 9732 23060 9738 23072
rect 9769 23069 9781 23072
rect 9815 23069 9827 23103
rect 9769 23063 9827 23069
rect 10410 23060 10416 23112
rect 10468 23060 10474 23112
rect 10962 23060 10968 23112
rect 11020 23100 11026 23112
rect 11057 23103 11115 23109
rect 11057 23100 11069 23103
rect 11020 23072 11069 23100
rect 11020 23060 11026 23072
rect 11057 23069 11069 23072
rect 11103 23069 11115 23103
rect 11057 23063 11115 23069
rect 7282 22992 7288 23044
rect 7340 22992 7346 23044
rect 7926 22992 7932 23044
rect 7984 22992 7990 23044
rect 11164 23032 11192 23140
rect 13173 23137 13185 23140
rect 13219 23137 13231 23171
rect 13173 23131 13231 23137
rect 13354 23128 13360 23180
rect 13412 23168 13418 23180
rect 16209 23171 16267 23177
rect 16209 23168 16221 23171
rect 13412 23140 16221 23168
rect 13412 23128 13418 23140
rect 16209 23137 16221 23140
rect 16255 23137 16267 23171
rect 18800 23168 18828 23199
rect 16209 23131 16267 23137
rect 16684 23140 18828 23168
rect 12894 23060 12900 23112
rect 12952 23100 12958 23112
rect 13449 23103 13507 23109
rect 13449 23100 13461 23103
rect 12952 23072 13461 23100
rect 12952 23060 12958 23072
rect 13449 23069 13461 23072
rect 13495 23069 13507 23103
rect 13449 23063 13507 23069
rect 13538 23060 13544 23112
rect 13596 23100 13602 23112
rect 13725 23103 13783 23109
rect 13725 23100 13737 23103
rect 13596 23072 13737 23100
rect 13596 23060 13602 23072
rect 13725 23069 13737 23072
rect 13771 23069 13783 23103
rect 13725 23063 13783 23069
rect 15102 23060 15108 23112
rect 15160 23060 15166 23112
rect 15562 23060 15568 23112
rect 15620 23060 15626 23112
rect 15654 23060 15660 23112
rect 15712 23100 15718 23112
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15712 23072 16037 23100
rect 15712 23060 15718 23072
rect 16025 23069 16037 23072
rect 16071 23100 16083 23103
rect 16684 23100 16712 23140
rect 16071 23072 16712 23100
rect 16071 23069 16083 23072
rect 16025 23063 16083 23069
rect 17402 23060 17408 23112
rect 17460 23100 17466 23112
rect 17957 23103 18015 23109
rect 17957 23100 17969 23103
rect 17460 23072 17969 23100
rect 17460 23060 17466 23072
rect 17957 23069 17969 23072
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 18966 23060 18972 23112
rect 19024 23060 19030 23112
rect 19426 23060 19432 23112
rect 19484 23060 19490 23112
rect 10980 23004 11192 23032
rect 10980 22976 11008 23004
rect 11882 22992 11888 23044
rect 11940 22992 11946 23044
rect 12437 23035 12495 23041
rect 12437 23001 12449 23035
rect 12483 23032 12495 23035
rect 12802 23032 12808 23044
rect 12483 23004 12808 23032
rect 12483 23001 12495 23004
rect 12437 22995 12495 23001
rect 12802 22992 12808 23004
rect 12860 22992 12866 23044
rect 12989 23035 13047 23041
rect 12989 23001 13001 23035
rect 13035 23032 13047 23035
rect 13035 23004 13676 23032
rect 13035 23001 13047 23004
rect 12989 22995 13047 23001
rect 13648 22976 13676 23004
rect 13998 22992 14004 23044
rect 14056 23032 14062 23044
rect 14369 23035 14427 23041
rect 14369 23032 14381 23035
rect 14056 23004 14381 23032
rect 14056 22992 14062 23004
rect 14369 23001 14381 23004
rect 14415 23001 14427 23035
rect 14369 22995 14427 23001
rect 16758 22992 16764 23044
rect 16816 22992 16822 23044
rect 17310 22992 17316 23044
rect 17368 22992 17374 23044
rect 18046 22992 18052 23044
rect 18104 23032 18110 23044
rect 18233 23035 18291 23041
rect 18233 23032 18245 23035
rect 18104 23004 18245 23032
rect 18104 22992 18110 23004
rect 18233 23001 18245 23004
rect 18279 23001 18291 23035
rect 18233 22995 18291 23001
rect 4614 22924 4620 22976
rect 4672 22924 4678 22976
rect 5442 22924 5448 22976
rect 5500 22924 5506 22976
rect 6733 22967 6791 22973
rect 6733 22933 6745 22967
rect 6779 22964 6791 22967
rect 7742 22964 7748 22976
rect 6779 22936 7748 22964
rect 6779 22933 6791 22936
rect 6733 22927 6791 22933
rect 7742 22924 7748 22936
rect 7800 22924 7806 22976
rect 8386 22924 8392 22976
rect 8444 22964 8450 22976
rect 8481 22967 8539 22973
rect 8481 22964 8493 22967
rect 8444 22936 8493 22964
rect 8444 22924 8450 22936
rect 8481 22933 8493 22936
rect 8527 22933 8539 22967
rect 8481 22927 8539 22933
rect 9950 22924 9956 22976
rect 10008 22924 10014 22976
rect 10597 22967 10655 22973
rect 10597 22933 10609 22967
rect 10643 22964 10655 22967
rect 10870 22964 10876 22976
rect 10643 22936 10876 22964
rect 10643 22933 10655 22936
rect 10597 22927 10655 22933
rect 10870 22924 10876 22936
rect 10928 22924 10934 22976
rect 10962 22924 10968 22976
rect 11020 22924 11026 22976
rect 11241 22967 11299 22973
rect 11241 22933 11253 22967
rect 11287 22964 11299 22967
rect 11698 22964 11704 22976
rect 11287 22936 11704 22964
rect 11287 22933 11299 22936
rect 11241 22927 11299 22933
rect 11698 22924 11704 22936
rect 11756 22924 11762 22976
rect 12618 22924 12624 22976
rect 12676 22924 12682 22976
rect 13078 22924 13084 22976
rect 13136 22924 13142 22976
rect 13630 22924 13636 22976
rect 13688 22924 13694 22976
rect 13906 22924 13912 22976
rect 13964 22924 13970 22976
rect 14550 22924 14556 22976
rect 14608 22964 14614 22976
rect 14921 22967 14979 22973
rect 14921 22964 14933 22967
rect 14608 22936 14933 22964
rect 14608 22924 14614 22936
rect 14921 22933 14933 22936
rect 14967 22933 14979 22967
rect 14921 22927 14979 22933
rect 15378 22924 15384 22976
rect 15436 22924 15442 22976
rect 15657 22967 15715 22973
rect 15657 22933 15669 22967
rect 15703 22964 15715 22967
rect 15746 22964 15752 22976
rect 15703 22936 15752 22964
rect 15703 22933 15715 22936
rect 15657 22927 15715 22933
rect 15746 22924 15752 22936
rect 15804 22924 15810 22976
rect 16114 22924 16120 22976
rect 16172 22924 16178 22976
rect 16482 22924 16488 22976
rect 16540 22964 16546 22976
rect 17773 22967 17831 22973
rect 17773 22964 17785 22967
rect 16540 22936 17785 22964
rect 16540 22924 16546 22936
rect 17773 22933 17785 22936
rect 17819 22933 17831 22967
rect 17773 22927 17831 22933
rect 19426 22924 19432 22976
rect 19484 22964 19490 22976
rect 19613 22967 19671 22973
rect 19613 22964 19625 22967
rect 19484 22936 19625 22964
rect 19484 22924 19490 22936
rect 19613 22933 19625 22936
rect 19659 22933 19671 22967
rect 19613 22927 19671 22933
rect 1104 22874 22356 22896
rect 1104 22822 4266 22874
rect 4318 22822 4330 22874
rect 4382 22822 4394 22874
rect 4446 22822 4458 22874
rect 4510 22822 4522 22874
rect 4574 22822 9579 22874
rect 9631 22822 9643 22874
rect 9695 22822 9707 22874
rect 9759 22822 9771 22874
rect 9823 22822 9835 22874
rect 9887 22822 14892 22874
rect 14944 22822 14956 22874
rect 15008 22822 15020 22874
rect 15072 22822 15084 22874
rect 15136 22822 15148 22874
rect 15200 22822 20205 22874
rect 20257 22822 20269 22874
rect 20321 22822 20333 22874
rect 20385 22822 20397 22874
rect 20449 22822 20461 22874
rect 20513 22822 22356 22874
rect 1104 22800 22356 22822
rect 7742 22720 7748 22772
rect 7800 22760 7806 22772
rect 7800 22732 8708 22760
rect 7800 22720 7806 22732
rect 7837 22695 7895 22701
rect 7837 22661 7849 22695
rect 7883 22692 7895 22695
rect 8527 22695 8585 22701
rect 8527 22692 8539 22695
rect 7883 22664 8539 22692
rect 7883 22661 7895 22664
rect 7837 22655 7895 22661
rect 8527 22661 8539 22664
rect 8573 22661 8585 22695
rect 8527 22655 8585 22661
rect 842 22584 848 22636
rect 900 22624 906 22636
rect 8386 22633 8392 22636
rect 1489 22627 1547 22633
rect 1489 22624 1501 22627
rect 900 22596 1501 22624
rect 900 22584 906 22596
rect 1489 22593 1501 22596
rect 1535 22593 1547 22627
rect 1489 22587 1547 22593
rect 8354 22627 8392 22633
rect 8354 22593 8366 22627
rect 8354 22587 8392 22593
rect 8386 22584 8392 22587
rect 8444 22584 8450 22636
rect 8680 22633 8708 22732
rect 13078 22720 13084 22772
rect 13136 22760 13142 22772
rect 13587 22763 13645 22769
rect 13587 22760 13599 22763
rect 13136 22732 13599 22760
rect 13136 22720 13142 22732
rect 13587 22729 13599 22732
rect 13633 22729 13645 22763
rect 13587 22723 13645 22729
rect 15335 22763 15393 22769
rect 15335 22729 15347 22763
rect 15381 22760 15393 22763
rect 16114 22760 16120 22772
rect 15381 22732 16120 22760
rect 15381 22729 15393 22732
rect 15335 22723 15393 22729
rect 16114 22720 16120 22732
rect 16172 22720 16178 22772
rect 13173 22695 13231 22701
rect 13173 22661 13185 22695
rect 13219 22692 13231 22695
rect 14090 22692 14096 22704
rect 13219 22664 14096 22692
rect 13219 22661 13231 22664
rect 13173 22655 13231 22661
rect 14090 22652 14096 22664
rect 14148 22652 14154 22704
rect 15841 22695 15899 22701
rect 15841 22661 15853 22695
rect 15887 22692 15899 22695
rect 15887 22664 16528 22692
rect 15887 22661 15899 22664
rect 15841 22655 15899 22661
rect 16500 22636 16528 22664
rect 8630 22627 8708 22633
rect 8630 22593 8642 22627
rect 8676 22596 8708 22627
rect 13081 22627 13139 22633
rect 8676 22593 8688 22596
rect 8630 22587 8688 22593
rect 13081 22593 13093 22627
rect 13127 22624 13139 22627
rect 13127 22596 13584 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 2041 22559 2099 22565
rect 2041 22525 2053 22559
rect 2087 22556 2099 22559
rect 2682 22556 2688 22568
rect 2087 22528 2688 22556
rect 2087 22525 2099 22528
rect 2041 22519 2099 22525
rect 2682 22516 2688 22528
rect 2740 22516 2746 22568
rect 7006 22516 7012 22568
rect 7064 22556 7070 22568
rect 8021 22559 8079 22565
rect 8021 22556 8033 22559
rect 7064 22528 8033 22556
rect 7064 22516 7070 22528
rect 8021 22525 8033 22528
rect 8067 22556 8079 22559
rect 10962 22556 10968 22568
rect 8067 22528 10968 22556
rect 8067 22525 8079 22528
rect 8021 22519 8079 22525
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 13354 22516 13360 22568
rect 13412 22516 13418 22568
rect 13556 22556 13584 22596
rect 13630 22584 13636 22636
rect 13688 22633 13694 22636
rect 13688 22627 13716 22633
rect 13704 22593 13716 22627
rect 13688 22587 13716 22593
rect 15264 22627 15322 22633
rect 15264 22593 15276 22627
rect 15310 22624 15322 22627
rect 15654 22624 15660 22636
rect 15310 22596 15660 22624
rect 15310 22593 15322 22596
rect 15264 22587 15322 22593
rect 13688 22584 13694 22587
rect 15654 22584 15660 22596
rect 15712 22584 15718 22636
rect 16482 22633 16488 22636
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22624 15991 22627
rect 16347 22627 16405 22633
rect 16347 22624 16359 22627
rect 15979 22596 16359 22624
rect 15979 22593 15991 22596
rect 15933 22587 15991 22593
rect 16347 22593 16359 22596
rect 16393 22593 16405 22627
rect 16347 22587 16405 22593
rect 16450 22627 16488 22633
rect 16450 22593 16462 22627
rect 16450 22587 16488 22593
rect 16482 22584 16488 22587
rect 16540 22584 16546 22636
rect 16666 22584 16672 22636
rect 16724 22584 16730 22636
rect 13906 22556 13912 22568
rect 13556 22528 13912 22556
rect 13906 22516 13912 22528
rect 13964 22516 13970 22568
rect 16071 22559 16129 22565
rect 16071 22525 16083 22559
rect 16117 22556 16129 22559
rect 16117 22528 16896 22556
rect 16117 22525 16129 22528
rect 16071 22519 16129 22525
rect 4890 22448 4896 22500
rect 4948 22488 4954 22500
rect 4948 22460 15608 22488
rect 4948 22448 4954 22460
rect 7098 22380 7104 22432
rect 7156 22420 7162 22432
rect 8294 22429 8300 22432
rect 7377 22423 7435 22429
rect 7377 22420 7389 22423
rect 7156 22392 7389 22420
rect 7156 22380 7162 22392
rect 7377 22389 7389 22392
rect 7423 22389 7435 22423
rect 7377 22383 7435 22389
rect 8251 22423 8300 22429
rect 8251 22389 8263 22423
rect 8297 22389 8300 22423
rect 8251 22383 8300 22389
rect 8294 22380 8300 22383
rect 8352 22380 8358 22432
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12713 22423 12771 22429
rect 12713 22420 12725 22423
rect 12492 22392 12725 22420
rect 12492 22380 12498 22392
rect 12713 22389 12725 22392
rect 12759 22389 12771 22423
rect 12713 22383 12771 22389
rect 15470 22380 15476 22432
rect 15528 22380 15534 22432
rect 15580 22420 15608 22460
rect 16666 22420 16672 22432
rect 15580 22392 16672 22420
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 16868 22429 16896 22528
rect 16853 22423 16911 22429
rect 16853 22389 16865 22423
rect 16899 22420 16911 22423
rect 19886 22420 19892 22432
rect 16899 22392 19892 22420
rect 16899 22389 16911 22392
rect 16853 22383 16911 22389
rect 19886 22380 19892 22392
rect 19944 22380 19950 22432
rect 1104 22330 22356 22352
rect 1104 22278 3606 22330
rect 3658 22278 3670 22330
rect 3722 22278 3734 22330
rect 3786 22278 3798 22330
rect 3850 22278 3862 22330
rect 3914 22278 8919 22330
rect 8971 22278 8983 22330
rect 9035 22278 9047 22330
rect 9099 22278 9111 22330
rect 9163 22278 9175 22330
rect 9227 22278 14232 22330
rect 14284 22278 14296 22330
rect 14348 22278 14360 22330
rect 14412 22278 14424 22330
rect 14476 22278 14488 22330
rect 14540 22278 19545 22330
rect 19597 22278 19609 22330
rect 19661 22278 19673 22330
rect 19725 22278 19737 22330
rect 19789 22278 19801 22330
rect 19853 22278 22356 22330
rect 1104 22256 22356 22278
rect 7098 22148 7104 22160
rect 6932 22120 7104 22148
rect 842 21972 848 22024
rect 900 22012 906 22024
rect 6932 22021 6960 22120
rect 7098 22108 7104 22120
rect 7156 22148 7162 22160
rect 7156 22120 8064 22148
rect 7156 22108 7162 22120
rect 7742 22040 7748 22092
rect 7800 22080 7806 22092
rect 7929 22083 7987 22089
rect 7929 22080 7941 22083
rect 7800 22052 7941 22080
rect 7800 22040 7806 22052
rect 7929 22049 7941 22052
rect 7975 22049 7987 22083
rect 8036 22080 8064 22120
rect 12618 22108 12624 22160
rect 12676 22148 12682 22160
rect 13541 22151 13599 22157
rect 13541 22148 13553 22151
rect 12676 22120 13553 22148
rect 12676 22108 12682 22120
rect 13541 22117 13553 22120
rect 13587 22117 13599 22151
rect 15746 22148 15752 22160
rect 13541 22111 13599 22117
rect 14844 22120 15752 22148
rect 8570 22080 8576 22092
rect 8036 22052 8576 22080
rect 7929 22043 7987 22049
rect 8570 22040 8576 22052
rect 8628 22040 8634 22092
rect 13262 22040 13268 22092
rect 13320 22040 13326 22092
rect 13906 22040 13912 22092
rect 13964 22040 13970 22092
rect 14090 22040 14096 22092
rect 14148 22089 14154 22092
rect 14148 22083 14197 22089
rect 14148 22049 14151 22083
rect 14185 22049 14197 22083
rect 14148 22043 14197 22049
rect 14737 22083 14795 22089
rect 14737 22049 14749 22083
rect 14783 22080 14795 22083
rect 14844 22080 14872 22120
rect 15746 22108 15752 22120
rect 15804 22148 15810 22160
rect 15804 22120 16160 22148
rect 15804 22108 15810 22120
rect 16132 22092 16160 22120
rect 14783 22052 14872 22080
rect 14921 22083 14979 22089
rect 14783 22049 14795 22052
rect 14737 22043 14795 22049
rect 14921 22049 14933 22083
rect 14967 22080 14979 22083
rect 15470 22080 15476 22092
rect 14967 22052 15476 22080
rect 14967 22049 14979 22052
rect 14921 22043 14979 22049
rect 14148 22040 14154 22043
rect 15470 22040 15476 22052
rect 15528 22040 15534 22092
rect 15562 22040 15568 22092
rect 15620 22040 15626 22092
rect 15654 22040 15660 22092
rect 15712 22080 15718 22092
rect 15841 22083 15899 22089
rect 15841 22080 15853 22083
rect 15712 22052 15853 22080
rect 15712 22040 15718 22052
rect 15841 22049 15853 22052
rect 15887 22049 15899 22083
rect 15841 22043 15899 22049
rect 16114 22040 16120 22092
rect 16172 22040 16178 22092
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 900 21984 1409 22012
rect 900 21972 906 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 6917 22015 6975 22021
rect 6917 21981 6929 22015
rect 6963 21981 6975 22015
rect 6917 21975 6975 21981
rect 7285 22015 7343 22021
rect 7285 21981 7297 22015
rect 7331 22012 7343 22015
rect 7837 22015 7895 22021
rect 7837 22012 7849 22015
rect 7331 21984 7849 22012
rect 7331 21981 7343 21984
rect 7285 21975 7343 21981
rect 7837 21981 7849 21984
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 8389 22015 8447 22021
rect 8389 21981 8401 22015
rect 8435 22012 8447 22015
rect 8478 22012 8484 22024
rect 8435 21984 8484 22012
rect 8435 21981 8447 21984
rect 8389 21975 8447 21981
rect 7101 21947 7159 21953
rect 7101 21913 7113 21947
rect 7147 21944 7159 21947
rect 7745 21947 7803 21953
rect 7147 21916 7696 21944
rect 7147 21913 7159 21916
rect 7101 21907 7159 21913
rect 1578 21836 1584 21888
rect 1636 21836 1642 21888
rect 7374 21836 7380 21888
rect 7432 21836 7438 21888
rect 7668 21876 7696 21916
rect 7745 21913 7757 21947
rect 7791 21944 7803 21947
rect 8205 21947 8263 21953
rect 8205 21944 8217 21947
rect 7791 21916 8217 21944
rect 7791 21913 7803 21916
rect 7745 21907 7803 21913
rect 8205 21913 8217 21916
rect 8251 21913 8263 21947
rect 8205 21907 8263 21913
rect 8404 21876 8432 21975
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 12253 22015 12311 22021
rect 12253 21981 12265 22015
rect 12299 22012 12311 22015
rect 13173 22015 13231 22021
rect 13173 22012 13185 22015
rect 12299 21984 13185 22012
rect 12299 21981 12311 21984
rect 12253 21975 12311 21981
rect 13173 21981 13185 21984
rect 13219 21981 13231 22015
rect 13173 21975 13231 21981
rect 13722 21972 13728 22024
rect 13780 21972 13786 22024
rect 13924 22012 13952 22040
rect 14226 22015 14284 22021
rect 14226 22012 14238 22015
rect 13924 21984 14238 22012
rect 14226 21981 14238 21984
rect 14272 21981 14284 22015
rect 15488 22012 15516 22040
rect 16209 22015 16267 22021
rect 16209 22012 16221 22015
rect 15488 21984 16221 22012
rect 14226 21975 14284 21981
rect 16209 21981 16221 21984
rect 16255 21981 16267 22015
rect 16209 21975 16267 21981
rect 12434 21904 12440 21956
rect 12492 21904 12498 21956
rect 12618 21904 12624 21956
rect 12676 21904 12682 21956
rect 13081 21947 13139 21953
rect 13081 21913 13093 21947
rect 13127 21944 13139 21947
rect 13909 21947 13967 21953
rect 13909 21944 13921 21947
rect 13127 21916 13921 21944
rect 13127 21913 13139 21916
rect 13081 21907 13139 21913
rect 13909 21913 13921 21916
rect 13955 21913 13967 21947
rect 13909 21907 13967 21913
rect 14553 21947 14611 21953
rect 14553 21913 14565 21947
rect 14599 21944 14611 21947
rect 15381 21947 15439 21953
rect 15381 21944 15393 21947
rect 14599 21916 15393 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 15381 21913 15393 21916
rect 15427 21913 15439 21947
rect 15381 21907 15439 21913
rect 7668 21848 8432 21876
rect 12710 21836 12716 21888
rect 12768 21836 12774 21888
rect 14642 21836 14648 21888
rect 14700 21876 14706 21888
rect 15013 21879 15071 21885
rect 15013 21876 15025 21879
rect 14700 21848 15025 21876
rect 14700 21836 14706 21848
rect 15013 21845 15025 21848
rect 15059 21845 15071 21879
rect 15013 21839 15071 21845
rect 15473 21879 15531 21885
rect 15473 21845 15485 21879
rect 15519 21876 15531 21879
rect 15930 21876 15936 21888
rect 15519 21848 15936 21876
rect 15519 21845 15531 21848
rect 15473 21839 15531 21845
rect 15930 21836 15936 21848
rect 15988 21836 15994 21888
rect 1104 21786 22356 21808
rect 1104 21734 4266 21786
rect 4318 21734 4330 21786
rect 4382 21734 4394 21786
rect 4446 21734 4458 21786
rect 4510 21734 4522 21786
rect 4574 21734 9579 21786
rect 9631 21734 9643 21786
rect 9695 21734 9707 21786
rect 9759 21734 9771 21786
rect 9823 21734 9835 21786
rect 9887 21734 14892 21786
rect 14944 21734 14956 21786
rect 15008 21734 15020 21786
rect 15072 21734 15084 21786
rect 15136 21734 15148 21786
rect 15200 21734 20205 21786
rect 20257 21734 20269 21786
rect 20321 21734 20333 21786
rect 20385 21734 20397 21786
rect 20449 21734 20461 21786
rect 20513 21734 22356 21786
rect 1104 21712 22356 21734
rect 5169 21675 5227 21681
rect 5169 21641 5181 21675
rect 5215 21672 5227 21675
rect 5442 21672 5448 21684
rect 5215 21644 5448 21672
rect 5215 21641 5227 21644
rect 5169 21635 5227 21641
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 8021 21675 8079 21681
rect 8021 21641 8033 21675
rect 8067 21672 8079 21675
rect 8294 21672 8300 21684
rect 8067 21644 8300 21672
rect 8067 21641 8079 21644
rect 8021 21635 8079 21641
rect 8294 21632 8300 21644
rect 8352 21632 8358 21684
rect 15930 21632 15936 21684
rect 15988 21632 15994 21684
rect 5460 21604 5488 21632
rect 5460 21576 5856 21604
rect 842 21496 848 21548
rect 900 21536 906 21548
rect 1489 21539 1547 21545
rect 1489 21536 1501 21539
rect 900 21508 1501 21536
rect 900 21496 906 21508
rect 1489 21505 1501 21508
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 4490 21539 4548 21545
rect 4490 21505 4502 21539
rect 4536 21536 4548 21539
rect 4614 21536 4620 21548
rect 4536 21508 4620 21536
rect 4536 21505 4548 21508
rect 4490 21499 4548 21505
rect 4614 21496 4620 21508
rect 4672 21496 4678 21548
rect 5828 21545 5856 21576
rect 5261 21539 5319 21545
rect 5261 21505 5273 21539
rect 5307 21536 5319 21539
rect 5675 21539 5733 21545
rect 5675 21536 5687 21539
rect 5307 21508 5687 21536
rect 5307 21505 5319 21508
rect 5261 21499 5319 21505
rect 5675 21505 5687 21508
rect 5721 21505 5733 21539
rect 5675 21499 5733 21505
rect 5778 21539 5856 21545
rect 5778 21505 5790 21539
rect 5824 21508 5856 21539
rect 5920 21576 8156 21604
rect 5824 21505 5836 21508
rect 5778 21499 5836 21505
rect 4154 21428 4160 21480
rect 4212 21468 4218 21480
rect 5445 21471 5503 21477
rect 5445 21468 5457 21471
rect 4212 21440 5457 21468
rect 4212 21428 4218 21440
rect 5445 21437 5457 21440
rect 5491 21468 5503 21471
rect 5920 21468 5948 21576
rect 7098 21496 7104 21548
rect 7156 21496 7162 21548
rect 7929 21539 7987 21545
rect 7929 21505 7941 21539
rect 7975 21536 7987 21539
rect 8018 21536 8024 21548
rect 7975 21508 8024 21536
rect 7975 21505 7987 21508
rect 7929 21499 7987 21505
rect 8018 21496 8024 21508
rect 8076 21496 8082 21548
rect 8128 21477 8156 21576
rect 8220 21576 8524 21604
rect 5491 21440 5948 21468
rect 7193 21471 7251 21477
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 8113 21471 8171 21477
rect 7239 21440 7604 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 1673 21403 1731 21409
rect 1673 21369 1685 21403
rect 1719 21400 1731 21403
rect 4982 21400 4988 21412
rect 1719 21372 4988 21400
rect 1719 21369 1731 21372
rect 1673 21363 1731 21369
rect 4982 21360 4988 21372
rect 5040 21360 5046 21412
rect 4387 21335 4445 21341
rect 4387 21301 4399 21335
rect 4433 21332 4445 21335
rect 4522 21332 4528 21344
rect 4433 21304 4528 21332
rect 4433 21301 4445 21304
rect 4387 21295 4445 21301
rect 4522 21292 4528 21304
rect 4580 21292 4586 21344
rect 4801 21335 4859 21341
rect 4801 21301 4813 21335
rect 4847 21332 4859 21335
rect 5534 21332 5540 21344
rect 4847 21304 5540 21332
rect 4847 21301 4859 21304
rect 4801 21295 4859 21301
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 7190 21292 7196 21344
rect 7248 21332 7254 21344
rect 7576 21341 7604 21440
rect 8113 21437 8125 21471
rect 8159 21437 8171 21471
rect 8113 21431 8171 21437
rect 7469 21335 7527 21341
rect 7469 21332 7481 21335
rect 7248 21304 7481 21332
rect 7248 21292 7254 21304
rect 7469 21301 7481 21304
rect 7515 21301 7527 21335
rect 7469 21295 7527 21301
rect 7561 21335 7619 21341
rect 7561 21301 7573 21335
rect 7607 21332 7619 21335
rect 8220 21332 8248 21576
rect 8496 21548 8524 21576
rect 15470 21564 15476 21616
rect 15528 21604 15534 21616
rect 16301 21607 16359 21613
rect 16301 21604 16313 21607
rect 15528 21576 16313 21604
rect 15528 21564 15534 21576
rect 16301 21573 16313 21576
rect 16347 21573 16359 21607
rect 16301 21567 16359 21573
rect 8478 21496 8484 21548
rect 8536 21536 8542 21548
rect 8573 21539 8631 21545
rect 8573 21536 8585 21539
rect 8536 21508 8585 21536
rect 8536 21496 8542 21508
rect 8573 21505 8585 21508
rect 8619 21505 8631 21539
rect 8573 21499 8631 21505
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 12805 21539 12863 21545
rect 12805 21536 12817 21539
rect 12676 21508 12817 21536
rect 12676 21496 12682 21508
rect 12805 21505 12817 21508
rect 12851 21505 12863 21539
rect 12805 21499 12863 21505
rect 15657 21539 15715 21545
rect 15657 21505 15669 21539
rect 15703 21536 15715 21539
rect 16114 21536 16120 21548
rect 15703 21508 16120 21536
rect 15703 21505 15715 21508
rect 15657 21499 15715 21505
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 12434 21428 12440 21480
rect 12492 21468 12498 21480
rect 12713 21471 12771 21477
rect 12713 21468 12725 21471
rect 12492 21440 12725 21468
rect 12492 21428 12498 21440
rect 12713 21437 12725 21440
rect 12759 21468 12771 21471
rect 13449 21471 13507 21477
rect 13449 21468 13461 21471
rect 12759 21440 13461 21468
rect 12759 21437 12771 21440
rect 12713 21431 12771 21437
rect 13449 21437 13461 21440
rect 13495 21468 13507 21471
rect 13722 21468 13728 21480
rect 13495 21440 13728 21468
rect 13495 21437 13507 21440
rect 13449 21431 13507 21437
rect 13722 21428 13728 21440
rect 13780 21428 13786 21480
rect 15470 21428 15476 21480
rect 15528 21428 15534 21480
rect 8389 21403 8447 21409
rect 8389 21369 8401 21403
rect 8435 21400 8447 21403
rect 8570 21400 8576 21412
rect 8435 21372 8576 21400
rect 8435 21369 8447 21372
rect 8389 21363 8447 21369
rect 8570 21360 8576 21372
rect 8628 21360 8634 21412
rect 12618 21360 12624 21412
rect 12676 21400 12682 21412
rect 13265 21403 13323 21409
rect 13265 21400 13277 21403
rect 12676 21372 13277 21400
rect 12676 21360 12682 21372
rect 13265 21369 13277 21372
rect 13311 21369 13323 21403
rect 13265 21363 13323 21369
rect 7607 21304 8248 21332
rect 7607 21301 7619 21304
rect 7561 21295 7619 21301
rect 8294 21292 8300 21344
rect 8352 21332 8358 21344
rect 8757 21335 8815 21341
rect 8757 21332 8769 21335
rect 8352 21304 8769 21332
rect 8352 21292 8358 21304
rect 8757 21301 8769 21304
rect 8803 21301 8815 21335
rect 8757 21295 8815 21301
rect 13170 21292 13176 21344
rect 13228 21292 13234 21344
rect 13446 21292 13452 21344
rect 13504 21332 13510 21344
rect 13633 21335 13691 21341
rect 13633 21332 13645 21335
rect 13504 21304 13645 21332
rect 13504 21292 13510 21304
rect 13633 21301 13645 21304
rect 13679 21301 13691 21335
rect 13633 21295 13691 21301
rect 15838 21292 15844 21344
rect 15896 21292 15902 21344
rect 1104 21242 22356 21264
rect 1104 21190 3606 21242
rect 3658 21190 3670 21242
rect 3722 21190 3734 21242
rect 3786 21190 3798 21242
rect 3850 21190 3862 21242
rect 3914 21190 8919 21242
rect 8971 21190 8983 21242
rect 9035 21190 9047 21242
rect 9099 21190 9111 21242
rect 9163 21190 9175 21242
rect 9227 21190 14232 21242
rect 14284 21190 14296 21242
rect 14348 21190 14360 21242
rect 14412 21190 14424 21242
rect 14476 21190 14488 21242
rect 14540 21190 19545 21242
rect 19597 21190 19609 21242
rect 19661 21190 19673 21242
rect 19725 21190 19737 21242
rect 19789 21190 19801 21242
rect 19853 21190 22356 21242
rect 1104 21168 22356 21190
rect 2682 21020 2688 21072
rect 2740 21060 2746 21072
rect 4890 21060 4896 21072
rect 2740 21032 4896 21060
rect 2740 21020 2746 21032
rect 4890 21020 4896 21032
rect 4948 21020 4954 21072
rect 15197 21063 15255 21069
rect 15197 21029 15209 21063
rect 15243 21060 15255 21063
rect 15654 21060 15660 21072
rect 15243 21032 15660 21060
rect 15243 21029 15255 21032
rect 15197 21023 15255 21029
rect 15654 21020 15660 21032
rect 15712 21020 15718 21072
rect 4522 20952 4528 21004
rect 4580 20952 4586 21004
rect 4706 20952 4712 21004
rect 4764 20952 4770 21004
rect 6822 20992 6828 21004
rect 4816 20964 6828 20992
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 4816 20924 4844 20964
rect 6822 20952 6828 20964
rect 6880 20952 6886 21004
rect 7190 20952 7196 21004
rect 7248 20992 7254 21004
rect 7285 20995 7343 21001
rect 7285 20992 7297 20995
rect 7248 20964 7297 20992
rect 7248 20952 7254 20964
rect 7285 20961 7297 20964
rect 7331 20961 7343 20995
rect 7285 20955 7343 20961
rect 18601 20995 18659 21001
rect 18601 20961 18613 20995
rect 18647 20992 18659 20995
rect 18647 20964 19104 20992
rect 18647 20961 18659 20964
rect 18601 20955 18659 20961
rect 1719 20896 4844 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 4890 20884 4896 20936
rect 4948 20884 4954 20936
rect 7006 20924 7012 20936
rect 5184 20896 7012 20924
rect 4433 20859 4491 20865
rect 4433 20825 4445 20859
rect 4479 20856 4491 20859
rect 4614 20856 4620 20868
rect 4479 20828 4620 20856
rect 4479 20825 4491 20828
rect 4433 20819 4491 20825
rect 4614 20816 4620 20828
rect 4672 20816 4678 20868
rect 4706 20816 4712 20868
rect 4764 20856 4770 20868
rect 5184 20865 5212 20896
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 7466 20884 7472 20936
rect 7524 20884 7530 20936
rect 8294 20884 8300 20936
rect 8352 20884 8358 20936
rect 13446 20884 13452 20936
rect 13504 20884 13510 20936
rect 13817 20927 13875 20933
rect 13817 20893 13829 20927
rect 13863 20924 13875 20927
rect 15286 20924 15292 20936
rect 13863 20896 15292 20924
rect 13863 20893 13875 20896
rect 13817 20887 13875 20893
rect 15286 20884 15292 20896
rect 15344 20924 15350 20936
rect 15381 20927 15439 20933
rect 15381 20924 15393 20927
rect 15344 20896 15393 20924
rect 15344 20884 15350 20896
rect 15381 20893 15393 20896
rect 15427 20893 15439 20927
rect 15381 20887 15439 20893
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 16117 20927 16175 20933
rect 16117 20924 16129 20927
rect 15611 20896 16129 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 16117 20893 16129 20896
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20924 16359 20927
rect 17126 20924 17132 20936
rect 16347 20896 17132 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 17126 20884 17132 20896
rect 17184 20924 17190 20936
rect 17405 20927 17463 20933
rect 17405 20924 17417 20927
rect 17184 20896 17417 20924
rect 17184 20884 17190 20896
rect 17405 20893 17417 20896
rect 17451 20893 17463 20927
rect 17405 20887 17463 20893
rect 17494 20884 17500 20936
rect 17552 20884 17558 20936
rect 18322 20884 18328 20936
rect 18380 20924 18386 20936
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 18380 20896 18429 20924
rect 18380 20884 18386 20896
rect 18417 20893 18429 20896
rect 18463 20924 18475 20927
rect 18877 20927 18935 20933
rect 18877 20924 18889 20927
rect 18463 20896 18889 20924
rect 18463 20893 18475 20896
rect 18417 20887 18475 20893
rect 18877 20893 18889 20896
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 19076 20868 19104 20964
rect 19886 20952 19892 21004
rect 19944 20992 19950 21004
rect 20530 20992 20536 21004
rect 19944 20964 20536 20992
rect 19944 20952 19950 20964
rect 20530 20952 20536 20964
rect 20588 20952 20594 21004
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 19484 20896 19625 20924
rect 19484 20884 19490 20896
rect 19613 20893 19625 20896
rect 19659 20924 19671 20927
rect 20190 20927 20248 20933
rect 20190 20924 20202 20927
rect 19659 20896 20202 20924
rect 19659 20893 19671 20896
rect 19613 20887 19671 20893
rect 20190 20893 20202 20896
rect 20236 20893 20248 20927
rect 20190 20887 20248 20893
rect 22002 20884 22008 20936
rect 22060 20884 22066 20936
rect 5169 20859 5227 20865
rect 5169 20856 5181 20859
rect 4764 20828 5181 20856
rect 4764 20816 4770 20828
rect 5169 20825 5181 20828
rect 5215 20825 5227 20859
rect 5169 20819 5227 20825
rect 5534 20816 5540 20868
rect 5592 20856 5598 20868
rect 5629 20859 5687 20865
rect 5629 20856 5641 20859
rect 5592 20828 5641 20856
rect 5592 20816 5598 20828
rect 5629 20825 5641 20828
rect 5675 20825 5687 20859
rect 5629 20819 5687 20825
rect 5718 20816 5724 20868
rect 5776 20856 5782 20868
rect 5813 20859 5871 20865
rect 5813 20856 5825 20859
rect 5776 20828 5825 20856
rect 5776 20816 5782 20828
rect 5813 20825 5825 20828
rect 5859 20825 5871 20859
rect 5813 20819 5871 20825
rect 7653 20859 7711 20865
rect 7653 20825 7665 20859
rect 7699 20856 7711 20859
rect 8113 20859 8171 20865
rect 8113 20856 8125 20859
rect 7699 20828 8125 20856
rect 7699 20825 7711 20828
rect 7653 20819 7711 20825
rect 8113 20825 8125 20828
rect 8159 20825 8171 20859
rect 8113 20819 8171 20825
rect 13630 20816 13636 20868
rect 13688 20816 13694 20868
rect 15838 20816 15844 20868
rect 15896 20856 15902 20868
rect 15933 20859 15991 20865
rect 15933 20856 15945 20859
rect 15896 20828 15945 20856
rect 15896 20816 15902 20828
rect 15933 20825 15945 20828
rect 15979 20825 15991 20859
rect 15933 20819 15991 20825
rect 17957 20859 18015 20865
rect 17957 20825 17969 20859
rect 18003 20856 18015 20859
rect 18598 20856 18604 20868
rect 18003 20828 18604 20856
rect 18003 20825 18015 20828
rect 17957 20819 18015 20825
rect 18598 20816 18604 20828
rect 18656 20816 18662 20868
rect 19058 20816 19064 20868
rect 19116 20856 19122 20868
rect 19116 20828 19288 20856
rect 19116 20816 19122 20828
rect 1486 20748 1492 20800
rect 1544 20748 1550 20800
rect 3970 20748 3976 20800
rect 4028 20788 4034 20800
rect 4065 20791 4123 20797
rect 4065 20788 4077 20791
rect 4028 20760 4077 20788
rect 4028 20748 4034 20760
rect 4065 20757 4077 20760
rect 4111 20757 4123 20791
rect 4065 20751 4123 20757
rect 5442 20748 5448 20800
rect 5500 20748 5506 20800
rect 7929 20791 7987 20797
rect 7929 20757 7941 20791
rect 7975 20788 7987 20791
rect 9306 20788 9312 20800
rect 7975 20760 9312 20788
rect 7975 20757 7987 20760
rect 7929 20751 7987 20757
rect 9306 20748 9312 20760
rect 9364 20748 9370 20800
rect 18230 20748 18236 20800
rect 18288 20748 18294 20800
rect 18690 20748 18696 20800
rect 18748 20748 18754 20800
rect 19260 20797 19288 20828
rect 19245 20791 19303 20797
rect 19245 20757 19257 20791
rect 19291 20757 19303 20791
rect 19245 20751 19303 20757
rect 19705 20791 19763 20797
rect 19705 20757 19717 20791
rect 19751 20788 19763 20791
rect 20119 20791 20177 20797
rect 20119 20788 20131 20791
rect 19751 20760 20131 20788
rect 19751 20757 19763 20760
rect 19705 20751 19763 20757
rect 20119 20757 20131 20760
rect 20165 20757 20177 20791
rect 20119 20751 20177 20757
rect 21818 20748 21824 20800
rect 21876 20748 21882 20800
rect 1104 20698 22356 20720
rect 1104 20646 4266 20698
rect 4318 20646 4330 20698
rect 4382 20646 4394 20698
rect 4446 20646 4458 20698
rect 4510 20646 4522 20698
rect 4574 20646 9579 20698
rect 9631 20646 9643 20698
rect 9695 20646 9707 20698
rect 9759 20646 9771 20698
rect 9823 20646 9835 20698
rect 9887 20646 14892 20698
rect 14944 20646 14956 20698
rect 15008 20646 15020 20698
rect 15072 20646 15084 20698
rect 15136 20646 15148 20698
rect 15200 20646 20205 20698
rect 20257 20646 20269 20698
rect 20321 20646 20333 20698
rect 20385 20646 20397 20698
rect 20449 20646 20461 20698
rect 20513 20646 22356 20698
rect 1104 20624 22356 20646
rect 5261 20587 5319 20593
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 5442 20584 5448 20596
rect 5307 20556 5448 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 5442 20544 5448 20556
rect 5500 20544 5506 20596
rect 9950 20544 9956 20596
rect 10008 20584 10014 20596
rect 10781 20587 10839 20593
rect 10781 20584 10793 20587
rect 10008 20556 10793 20584
rect 10008 20544 10014 20556
rect 10781 20553 10793 20556
rect 10827 20553 10839 20587
rect 10781 20547 10839 20553
rect 4249 20519 4307 20525
rect 4249 20485 4261 20519
rect 4295 20516 4307 20519
rect 5813 20519 5871 20525
rect 5813 20516 5825 20519
rect 4295 20488 5825 20516
rect 4295 20485 4307 20488
rect 4249 20479 4307 20485
rect 5813 20485 5825 20488
rect 5859 20485 5871 20519
rect 10796 20516 10824 20547
rect 18230 20544 18236 20596
rect 18288 20584 18294 20596
rect 18325 20587 18383 20593
rect 18325 20584 18337 20587
rect 18288 20556 18337 20584
rect 18288 20544 18294 20556
rect 18325 20553 18337 20556
rect 18371 20553 18383 20587
rect 18325 20547 18383 20553
rect 18417 20587 18475 20593
rect 18417 20553 18429 20587
rect 18463 20584 18475 20587
rect 18690 20584 18696 20596
rect 18463 20556 18696 20584
rect 18463 20553 18475 20556
rect 18417 20547 18475 20553
rect 18690 20544 18696 20556
rect 18748 20544 18754 20596
rect 19245 20587 19303 20593
rect 19245 20584 19257 20587
rect 18984 20556 19257 20584
rect 10796 20488 11677 20516
rect 5813 20479 5871 20485
rect 3970 20448 3976 20460
rect 3896 20420 3976 20448
rect 3896 20389 3924 20420
rect 3970 20408 3976 20420
rect 4028 20448 4034 20460
rect 4525 20451 4583 20457
rect 4525 20448 4537 20451
rect 4028 20420 4537 20448
rect 4028 20408 4034 20420
rect 4525 20417 4537 20420
rect 4571 20448 4583 20451
rect 4571 20420 5304 20448
rect 4571 20417 4583 20420
rect 4525 20411 4583 20417
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20349 3939 20383
rect 3881 20343 3939 20349
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 4111 20352 4629 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 4617 20349 4629 20352
rect 4663 20380 4675 20383
rect 5169 20383 5227 20389
rect 4663 20352 5120 20380
rect 4663 20349 4675 20352
rect 4617 20343 4675 20349
rect 4798 20204 4804 20256
rect 4856 20244 4862 20256
rect 4893 20247 4951 20253
rect 4893 20244 4905 20247
rect 4856 20216 4905 20244
rect 4856 20204 4862 20216
rect 4893 20213 4905 20216
rect 4939 20213 4951 20247
rect 5092 20244 5120 20352
rect 5169 20349 5181 20383
rect 5215 20349 5227 20383
rect 5276 20380 5304 20420
rect 5350 20408 5356 20460
rect 5408 20408 5414 20460
rect 5994 20408 6000 20460
rect 6052 20408 6058 20460
rect 6181 20451 6239 20457
rect 6181 20417 6193 20451
rect 6227 20448 6239 20451
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 6227 20420 7297 20448
rect 6227 20417 6239 20420
rect 6181 20411 6239 20417
rect 7285 20417 7297 20420
rect 7331 20448 7343 20451
rect 7466 20448 7472 20460
rect 7331 20420 7472 20448
rect 7331 20417 7343 20420
rect 7285 20411 7343 20417
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 9306 20408 9312 20460
rect 9364 20408 9370 20460
rect 9398 20408 9404 20460
rect 9456 20408 9462 20460
rect 11649 20457 11677 20488
rect 13630 20476 13636 20528
rect 13688 20476 13694 20528
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20448 10931 20451
rect 11563 20451 11621 20457
rect 11563 20448 11575 20451
rect 10919 20420 11575 20448
rect 10919 20417 10931 20420
rect 10873 20411 10931 20417
rect 11563 20417 11575 20420
rect 11609 20417 11621 20451
rect 11649 20451 11708 20457
rect 11649 20420 11662 20451
rect 11563 20411 11621 20417
rect 11650 20417 11662 20420
rect 11696 20417 11708 20451
rect 11650 20411 11708 20417
rect 13170 20408 13176 20460
rect 13228 20408 13234 20460
rect 15286 20408 15292 20460
rect 15344 20408 15350 20460
rect 17126 20408 17132 20460
rect 17184 20408 17190 20460
rect 18322 20408 18328 20460
rect 18380 20448 18386 20460
rect 18984 20457 19012 20556
rect 19245 20553 19257 20556
rect 19291 20553 19303 20587
rect 19245 20547 19303 20553
rect 19613 20519 19671 20525
rect 19613 20485 19625 20519
rect 19659 20516 19671 20519
rect 19659 20488 20300 20516
rect 19659 20485 19671 20488
rect 19613 20479 19671 20485
rect 20272 20457 20300 20488
rect 18969 20451 19027 20457
rect 18969 20448 18981 20451
rect 18380 20420 18981 20448
rect 18380 20408 18386 20420
rect 18969 20417 18981 20420
rect 19015 20417 19027 20451
rect 18969 20411 19027 20417
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20448 19763 20451
rect 20119 20451 20177 20457
rect 20119 20448 20131 20451
rect 19751 20420 20131 20448
rect 19751 20417 19763 20420
rect 19705 20411 19763 20417
rect 20119 20417 20131 20420
rect 20165 20417 20177 20451
rect 20119 20411 20177 20417
rect 20222 20451 20300 20457
rect 20222 20417 20234 20451
rect 20268 20448 20300 20451
rect 21818 20448 21824 20460
rect 20268 20420 21824 20448
rect 20268 20417 20280 20420
rect 20222 20411 20280 20417
rect 21818 20408 21824 20420
rect 21876 20408 21882 20460
rect 5626 20380 5632 20392
rect 5276 20352 5632 20380
rect 5169 20343 5227 20349
rect 5184 20312 5212 20343
rect 5626 20340 5632 20352
rect 5684 20340 5690 20392
rect 7190 20340 7196 20392
rect 7248 20340 7254 20392
rect 9861 20383 9919 20389
rect 9861 20349 9873 20383
rect 9907 20380 9919 20383
rect 10778 20380 10784 20392
rect 9907 20352 10784 20380
rect 9907 20349 9919 20352
rect 9861 20343 9919 20349
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 10962 20340 10968 20392
rect 11020 20340 11026 20392
rect 13078 20340 13084 20392
rect 13136 20340 13142 20392
rect 15381 20383 15439 20389
rect 15381 20349 15393 20383
rect 15427 20380 15439 20383
rect 15654 20380 15660 20392
rect 15427 20352 15660 20380
rect 15427 20349 15439 20352
rect 15381 20343 15439 20349
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 17221 20383 17279 20389
rect 17221 20349 17233 20383
rect 17267 20380 17279 20383
rect 17494 20380 17500 20392
rect 17267 20352 17500 20380
rect 17267 20349 17279 20352
rect 17221 20343 17279 20349
rect 17494 20340 17500 20352
rect 17552 20380 17558 20392
rect 17862 20380 17868 20392
rect 17552 20352 17868 20380
rect 17552 20340 17558 20352
rect 17862 20340 17868 20352
rect 17920 20340 17926 20392
rect 18414 20340 18420 20392
rect 18472 20380 18478 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18472 20352 18521 20380
rect 18472 20340 18478 20352
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 18509 20343 18567 20349
rect 19889 20383 19947 20389
rect 19889 20349 19901 20383
rect 19935 20380 19947 20383
rect 20622 20380 20628 20392
rect 19935 20352 20628 20380
rect 19935 20349 19947 20352
rect 19889 20343 19947 20349
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 7834 20312 7840 20324
rect 5184 20284 7840 20312
rect 7834 20272 7840 20284
rect 7892 20272 7898 20324
rect 10686 20272 10692 20324
rect 10744 20312 10750 20324
rect 10980 20312 11008 20340
rect 10744 20284 11008 20312
rect 10744 20272 10750 20284
rect 18230 20272 18236 20324
rect 18288 20312 18294 20324
rect 19058 20312 19064 20324
rect 18288 20284 19064 20312
rect 18288 20272 18294 20284
rect 19058 20272 19064 20284
rect 19116 20312 19122 20324
rect 19153 20315 19211 20321
rect 19153 20312 19165 20315
rect 19116 20284 19165 20312
rect 19116 20272 19122 20284
rect 19153 20281 19165 20284
rect 19199 20281 19211 20315
rect 19153 20275 19211 20281
rect 5534 20244 5540 20256
rect 5092 20216 5540 20244
rect 4893 20207 4951 20213
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 5718 20204 5724 20256
rect 5776 20204 5782 20256
rect 7558 20204 7564 20256
rect 7616 20244 7622 20256
rect 7653 20247 7711 20253
rect 7653 20244 7665 20247
rect 7616 20216 7665 20244
rect 7616 20204 7622 20216
rect 7653 20213 7665 20216
rect 7699 20213 7711 20247
rect 7653 20207 7711 20213
rect 10410 20204 10416 20256
rect 10468 20204 10474 20256
rect 14921 20247 14979 20253
rect 14921 20213 14933 20247
rect 14967 20244 14979 20247
rect 15194 20244 15200 20256
rect 14967 20216 15200 20244
rect 14967 20213 14979 20216
rect 14921 20207 14979 20213
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 16758 20204 16764 20256
rect 16816 20204 16822 20256
rect 17034 20204 17040 20256
rect 17092 20244 17098 20256
rect 17957 20247 18015 20253
rect 17957 20244 17969 20247
rect 17092 20216 17969 20244
rect 17092 20204 17098 20216
rect 17957 20213 17969 20216
rect 18003 20213 18015 20247
rect 17957 20207 18015 20213
rect 18785 20247 18843 20253
rect 18785 20213 18797 20247
rect 18831 20244 18843 20247
rect 18874 20244 18880 20256
rect 18831 20216 18880 20244
rect 18831 20213 18843 20216
rect 18785 20207 18843 20213
rect 18874 20204 18880 20216
rect 18932 20204 18938 20256
rect 1104 20154 22356 20176
rect 1104 20102 3606 20154
rect 3658 20102 3670 20154
rect 3722 20102 3734 20154
rect 3786 20102 3798 20154
rect 3850 20102 3862 20154
rect 3914 20102 8919 20154
rect 8971 20102 8983 20154
rect 9035 20102 9047 20154
rect 9099 20102 9111 20154
rect 9163 20102 9175 20154
rect 9227 20102 14232 20154
rect 14284 20102 14296 20154
rect 14348 20102 14360 20154
rect 14412 20102 14424 20154
rect 14476 20102 14488 20154
rect 14540 20102 19545 20154
rect 19597 20102 19609 20154
rect 19661 20102 19673 20154
rect 19725 20102 19737 20154
rect 19789 20102 19801 20154
rect 19853 20102 22356 20154
rect 1104 20080 22356 20102
rect 5261 20043 5319 20049
rect 5261 20009 5273 20043
rect 5307 20040 5319 20043
rect 5994 20040 6000 20052
rect 5307 20012 6000 20040
rect 5307 20009 5319 20012
rect 5261 20003 5319 20009
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 13354 20040 13360 20052
rect 12176 20012 13360 20040
rect 5350 19932 5356 19984
rect 5408 19972 5414 19984
rect 10689 19975 10747 19981
rect 5408 19944 6040 19972
rect 5408 19932 5414 19944
rect 4798 19864 4804 19916
rect 4856 19904 4862 19916
rect 4856 19876 5120 19904
rect 4856 19864 4862 19876
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 1719 19808 2774 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 2746 19768 2774 19808
rect 4982 19796 4988 19848
rect 5040 19796 5046 19848
rect 5092 19845 5120 19876
rect 5626 19864 5632 19916
rect 5684 19864 5690 19916
rect 6012 19913 6040 19944
rect 10689 19941 10701 19975
rect 10735 19972 10747 19975
rect 10735 19944 10824 19972
rect 10735 19941 10747 19944
rect 10689 19935 10747 19941
rect 5997 19907 6055 19913
rect 5997 19873 6009 19907
rect 6043 19873 6055 19907
rect 5997 19867 6055 19873
rect 7834 19864 7840 19916
rect 7892 19864 7898 19916
rect 8754 19864 8760 19916
rect 8812 19904 8818 19916
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 8812 19876 8953 19904
rect 8812 19864 8818 19876
rect 8941 19873 8953 19876
rect 8987 19873 8999 19907
rect 8941 19867 8999 19873
rect 9398 19864 9404 19916
rect 9456 19904 9462 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9456 19876 9689 19904
rect 9456 19864 9462 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19904 10195 19907
rect 10226 19904 10232 19916
rect 10183 19876 10232 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 10226 19864 10232 19876
rect 10284 19904 10290 19916
rect 10796 19904 10824 19944
rect 10284 19876 10824 19904
rect 10284 19864 10290 19876
rect 5077 19839 5135 19845
rect 5077 19805 5089 19839
rect 5123 19805 5135 19839
rect 5077 19799 5135 19805
rect 5534 19796 5540 19848
rect 5592 19836 5598 19848
rect 5813 19839 5871 19845
rect 5813 19836 5825 19839
rect 5592 19808 5825 19836
rect 5592 19796 5598 19808
rect 5813 19805 5825 19808
rect 5859 19805 5871 19839
rect 5813 19799 5871 19805
rect 7558 19796 7564 19848
rect 7616 19796 7622 19848
rect 7653 19839 7711 19845
rect 7653 19805 7665 19839
rect 7699 19836 7711 19839
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 7699 19808 8033 19836
rect 7699 19805 7711 19808
rect 7653 19799 7711 19805
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 9306 19796 9312 19848
rect 9364 19796 9370 19848
rect 10042 19796 10048 19848
rect 10100 19836 10106 19848
rect 10796 19836 10824 19876
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19904 11391 19907
rect 12176 19904 12204 20012
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 15562 20000 15568 20052
rect 15620 20040 15626 20052
rect 15841 20043 15899 20049
rect 15841 20040 15853 20043
rect 15620 20012 15853 20040
rect 15620 20000 15626 20012
rect 15841 20009 15853 20012
rect 15887 20040 15899 20043
rect 15887 20012 16574 20040
rect 15887 20009 15899 20012
rect 15841 20003 15899 20009
rect 12805 19975 12863 19981
rect 12805 19941 12817 19975
rect 12851 19972 12863 19975
rect 13814 19972 13820 19984
rect 12851 19944 13820 19972
rect 12851 19941 12863 19944
rect 12805 19935 12863 19941
rect 13814 19932 13820 19944
rect 13872 19932 13878 19984
rect 11379 19876 12204 19904
rect 12253 19907 12311 19913
rect 11379 19873 11391 19876
rect 11333 19867 11391 19873
rect 12253 19873 12265 19907
rect 12299 19904 12311 19907
rect 12526 19904 12532 19916
rect 12299 19876 12532 19904
rect 12299 19873 12311 19876
rect 12253 19867 12311 19873
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 13262 19864 13268 19916
rect 13320 19904 13326 19916
rect 13446 19904 13452 19916
rect 13320 19876 13452 19904
rect 13320 19864 13326 19876
rect 13446 19864 13452 19876
rect 13504 19864 13510 19916
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19904 15531 19907
rect 15580 19904 15608 20000
rect 16546 19972 16574 20012
rect 17862 20000 17868 20052
rect 17920 20000 17926 20052
rect 18414 19972 18420 19984
rect 16546 19944 18420 19972
rect 16592 19913 16620 19944
rect 18414 19932 18420 19944
rect 18472 19932 18478 19984
rect 15519 19876 15608 19904
rect 16577 19907 16635 19913
rect 15519 19873 15531 19876
rect 15473 19867 15531 19873
rect 16577 19873 16589 19907
rect 16623 19904 16635 19907
rect 17221 19907 17279 19913
rect 16623 19876 16657 19904
rect 16623 19873 16635 19876
rect 16577 19867 16635 19873
rect 17221 19873 17233 19907
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 12437 19839 12495 19845
rect 10100 19808 10456 19836
rect 10796 19808 11744 19836
rect 10100 19796 10106 19808
rect 10428 19780 10456 19808
rect 7006 19768 7012 19780
rect 2746 19740 7012 19768
rect 7006 19728 7012 19740
rect 7064 19728 7070 19780
rect 10410 19728 10416 19780
rect 10468 19768 10474 19780
rect 11716 19777 11744 19808
rect 12437 19805 12449 19839
rect 12483 19836 12495 19839
rect 12710 19836 12716 19848
rect 12483 19808 12716 19836
rect 12483 19805 12495 19808
rect 12437 19799 12495 19805
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 13725 19839 13783 19845
rect 13725 19836 13737 19839
rect 13403 19808 13737 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 13725 19805 13737 19808
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 14090 19796 14096 19848
rect 14148 19836 14154 19848
rect 14645 19839 14703 19845
rect 14645 19836 14657 19839
rect 14148 19808 14657 19836
rect 14148 19796 14154 19808
rect 14645 19805 14657 19808
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 15194 19796 15200 19848
rect 15252 19796 15258 19848
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19836 15347 19839
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 15335 19808 16037 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 16025 19805 16037 19808
rect 16071 19805 16083 19839
rect 16025 19799 16083 19805
rect 16758 19796 16764 19848
rect 16816 19796 16822 19848
rect 11517 19771 11575 19777
rect 11517 19768 11529 19771
rect 10468 19740 11529 19768
rect 10468 19728 10474 19740
rect 11517 19737 11529 19740
rect 11563 19737 11575 19771
rect 11517 19731 11575 19737
rect 11701 19771 11759 19777
rect 11701 19737 11713 19771
rect 11747 19737 11759 19771
rect 11701 19731 11759 19737
rect 12345 19771 12403 19777
rect 12345 19737 12357 19771
rect 12391 19768 12403 19771
rect 12391 19740 12940 19768
rect 12391 19737 12403 19740
rect 12345 19731 12403 19737
rect 842 19660 848 19712
rect 900 19700 906 19712
rect 1489 19703 1547 19709
rect 1489 19700 1501 19703
rect 900 19672 1501 19700
rect 900 19660 906 19672
rect 1489 19669 1501 19672
rect 1535 19669 1547 19703
rect 1489 19663 1547 19669
rect 7193 19703 7251 19709
rect 7193 19669 7205 19703
rect 7239 19700 7251 19703
rect 7282 19700 7288 19712
rect 7239 19672 7288 19700
rect 7239 19669 7251 19672
rect 7193 19663 7251 19669
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 11054 19660 11060 19712
rect 11112 19660 11118 19712
rect 11146 19660 11152 19712
rect 11204 19660 11210 19712
rect 11238 19660 11244 19712
rect 11296 19700 11302 19712
rect 12912 19709 12940 19740
rect 14458 19728 14464 19780
rect 14516 19728 14522 19780
rect 15470 19728 15476 19780
rect 15528 19768 15534 19780
rect 15749 19771 15807 19777
rect 15749 19768 15761 19771
rect 15528 19740 15761 19768
rect 15528 19728 15534 19740
rect 15749 19737 15761 19740
rect 15795 19737 15807 19771
rect 15749 19731 15807 19737
rect 16669 19771 16727 19777
rect 16669 19737 16681 19771
rect 16715 19768 16727 19771
rect 17236 19768 17264 19867
rect 18322 19864 18328 19916
rect 18380 19864 18386 19916
rect 18230 19796 18236 19848
rect 18288 19796 18294 19848
rect 18598 19796 18604 19848
rect 18656 19836 18662 19848
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 18656 19808 18705 19836
rect 18656 19796 18662 19808
rect 18693 19805 18705 19808
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 18874 19796 18880 19848
rect 18932 19796 18938 19848
rect 22002 19796 22008 19848
rect 22060 19796 22066 19848
rect 16715 19740 17264 19768
rect 16715 19737 16727 19740
rect 16669 19731 16727 19737
rect 11885 19703 11943 19709
rect 11885 19700 11897 19703
rect 11296 19672 11897 19700
rect 11296 19660 11302 19672
rect 11885 19669 11897 19672
rect 11931 19669 11943 19703
rect 11885 19663 11943 19669
rect 12897 19703 12955 19709
rect 12897 19669 12909 19703
rect 12943 19669 12955 19703
rect 12897 19663 12955 19669
rect 13262 19660 13268 19712
rect 13320 19660 13326 19712
rect 14734 19660 14740 19712
rect 14792 19700 14798 19712
rect 14829 19703 14887 19709
rect 14829 19700 14841 19703
rect 14792 19672 14841 19700
rect 14792 19660 14798 19672
rect 14829 19669 14841 19672
rect 14875 19669 14887 19703
rect 14829 19663 14887 19669
rect 17126 19660 17132 19712
rect 17184 19660 17190 19712
rect 18506 19660 18512 19712
rect 18564 19660 18570 19712
rect 21818 19660 21824 19712
rect 21876 19660 21882 19712
rect 1104 19610 22356 19632
rect 1104 19558 4266 19610
rect 4318 19558 4330 19610
rect 4382 19558 4394 19610
rect 4446 19558 4458 19610
rect 4510 19558 4522 19610
rect 4574 19558 9579 19610
rect 9631 19558 9643 19610
rect 9695 19558 9707 19610
rect 9759 19558 9771 19610
rect 9823 19558 9835 19610
rect 9887 19558 14892 19610
rect 14944 19558 14956 19610
rect 15008 19558 15020 19610
rect 15072 19558 15084 19610
rect 15136 19558 15148 19610
rect 15200 19558 20205 19610
rect 20257 19558 20269 19610
rect 20321 19558 20333 19610
rect 20385 19558 20397 19610
rect 20449 19558 20461 19610
rect 20513 19558 22356 19610
rect 1104 19536 22356 19558
rect 7282 19456 7288 19508
rect 7340 19456 7346 19508
rect 7374 19456 7380 19508
rect 7432 19456 7438 19508
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 10134 19456 10140 19508
rect 10192 19456 10198 19508
rect 10229 19499 10287 19505
rect 10229 19465 10241 19499
rect 10275 19496 10287 19499
rect 10275 19468 11100 19496
rect 10275 19465 10287 19468
rect 10229 19459 10287 19465
rect 7466 19428 7472 19440
rect 2746 19400 7472 19428
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 2746 19360 2774 19400
rect 7466 19388 7472 19400
rect 7524 19388 7530 19440
rect 9309 19431 9367 19437
rect 9309 19397 9321 19431
rect 9355 19428 9367 19431
rect 10597 19431 10655 19437
rect 10597 19428 10609 19431
rect 9355 19400 10609 19428
rect 9355 19397 9367 19400
rect 9309 19391 9367 19397
rect 10597 19397 10609 19400
rect 10643 19397 10655 19431
rect 10597 19391 10655 19397
rect 10778 19388 10784 19440
rect 10836 19388 10842 19440
rect 11072 19428 11100 19468
rect 11146 19456 11152 19508
rect 11204 19496 11210 19508
rect 11563 19499 11621 19505
rect 11563 19496 11575 19499
rect 11204 19468 11575 19496
rect 11204 19456 11210 19468
rect 11563 19465 11575 19468
rect 11609 19465 11621 19499
rect 11563 19459 11621 19465
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 13541 19499 13599 19505
rect 13541 19496 13553 19499
rect 12860 19468 13553 19496
rect 12860 19456 12866 19468
rect 13541 19465 13553 19468
rect 13587 19465 13599 19499
rect 13541 19459 13599 19465
rect 13814 19456 13820 19508
rect 13872 19456 13878 19508
rect 13998 19456 14004 19508
rect 14056 19456 14062 19508
rect 14277 19499 14335 19505
rect 14277 19465 14289 19499
rect 14323 19465 14335 19499
rect 14277 19459 14335 19465
rect 11238 19428 11244 19440
rect 11072 19400 11244 19428
rect 11238 19388 11244 19400
rect 11296 19388 11302 19440
rect 13832 19428 13860 19456
rect 13740 19400 13860 19428
rect 1719 19332 2774 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 4982 19320 4988 19372
rect 5040 19360 5046 19372
rect 5169 19363 5227 19369
rect 5169 19360 5181 19363
rect 5040 19332 5181 19360
rect 5040 19320 5046 19332
rect 5169 19329 5181 19332
rect 5215 19329 5227 19363
rect 8570 19360 8576 19372
rect 5169 19323 5227 19329
rect 8220 19332 8576 19360
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 4154 19292 4160 19304
rect 2924 19264 4160 19292
rect 2924 19252 2930 19264
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 4798 19252 4804 19304
rect 4856 19292 4862 19304
rect 5077 19295 5135 19301
rect 5077 19292 5089 19295
rect 4856 19264 5089 19292
rect 4856 19252 4862 19264
rect 5077 19261 5089 19264
rect 5123 19261 5135 19295
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 5077 19255 5135 19261
rect 6886 19264 7205 19292
rect 5810 19184 5816 19236
rect 5868 19224 5874 19236
rect 6886 19224 6914 19264
rect 7193 19261 7205 19264
rect 7239 19292 7251 19295
rect 8220 19292 8248 19332
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 9416 19332 10180 19360
rect 7239 19264 8248 19292
rect 8297 19295 8355 19301
rect 7239 19261 7251 19264
rect 7193 19255 7251 19261
rect 8297 19261 8309 19295
rect 8343 19292 8355 19295
rect 8849 19295 8907 19301
rect 8849 19292 8861 19295
rect 8343 19264 8861 19292
rect 8343 19261 8355 19264
rect 8297 19255 8355 19261
rect 8849 19261 8861 19264
rect 8895 19261 8907 19295
rect 8849 19255 8907 19261
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19292 9091 19295
rect 9416 19292 9444 19332
rect 9079 19264 9444 19292
rect 9493 19295 9551 19301
rect 9079 19261 9091 19264
rect 9033 19255 9091 19261
rect 9493 19261 9505 19295
rect 9539 19261 9551 19295
rect 9493 19255 9551 19261
rect 9677 19295 9735 19301
rect 9677 19261 9689 19295
rect 9723 19292 9735 19295
rect 10042 19292 10048 19304
rect 9723 19264 10048 19292
rect 9723 19261 9735 19264
rect 9677 19255 9735 19261
rect 5868 19196 6914 19224
rect 5868 19184 5874 19196
rect 7834 19184 7840 19236
rect 7892 19224 7898 19236
rect 9048 19224 9076 19255
rect 7892 19196 9076 19224
rect 9508 19224 9536 19255
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 10152 19292 10180 19332
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11634 19363 11692 19369
rect 11634 19360 11646 19363
rect 11112 19332 11646 19360
rect 11112 19320 11118 19332
rect 11634 19329 11646 19332
rect 11680 19329 11692 19363
rect 11634 19323 11692 19329
rect 13078 19320 13084 19372
rect 13136 19360 13142 19372
rect 13538 19360 13544 19372
rect 13136 19332 13544 19360
rect 13136 19320 13142 19332
rect 13538 19320 13544 19332
rect 13596 19320 13602 19372
rect 13740 19369 13768 19400
rect 13725 19363 13783 19369
rect 13725 19329 13737 19363
rect 13771 19329 13783 19363
rect 13725 19323 13783 19329
rect 13817 19363 13875 19369
rect 13817 19329 13829 19363
rect 13863 19360 13875 19363
rect 13906 19360 13912 19372
rect 13863 19332 13912 19360
rect 13863 19329 13875 19332
rect 13817 19323 13875 19329
rect 13906 19320 13912 19332
rect 13964 19360 13970 19372
rect 14292 19360 14320 19459
rect 14642 19456 14648 19508
rect 14700 19456 14706 19508
rect 14734 19456 14740 19508
rect 14792 19456 14798 19508
rect 15838 19456 15844 19508
rect 15896 19496 15902 19508
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 15896 19468 16681 19496
rect 15896 19456 15902 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 16669 19459 16727 19465
rect 17034 19456 17040 19508
rect 17092 19456 17098 19508
rect 17126 19456 17132 19508
rect 17184 19456 17190 19508
rect 21634 19456 21640 19508
rect 21692 19496 21698 19508
rect 21821 19499 21879 19505
rect 21821 19496 21833 19499
rect 21692 19468 21833 19496
rect 21692 19456 21698 19468
rect 21821 19465 21833 19468
rect 21867 19465 21879 19499
rect 21821 19459 21879 19465
rect 13964 19332 14320 19360
rect 13964 19320 13970 19332
rect 22002 19320 22008 19372
rect 22060 19320 22066 19372
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 10152 19264 10333 19292
rect 10321 19261 10333 19264
rect 10367 19261 10379 19295
rect 10321 19255 10379 19261
rect 13170 19252 13176 19304
rect 13228 19252 13234 19304
rect 13262 19252 13268 19304
rect 13320 19292 13326 19304
rect 13449 19295 13507 19301
rect 13449 19292 13461 19295
rect 13320 19264 13461 19292
rect 13320 19252 13326 19264
rect 13449 19261 13461 19264
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14516 19264 14933 19292
rect 14516 19252 14522 19264
rect 14921 19261 14933 19264
rect 14967 19292 14979 19295
rect 17313 19295 17371 19301
rect 17313 19292 17325 19295
rect 14967 19264 17325 19292
rect 14967 19261 14979 19264
rect 14921 19255 14979 19261
rect 17313 19261 17325 19264
rect 17359 19292 17371 19295
rect 17402 19292 17408 19304
rect 17359 19264 17408 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 10226 19224 10232 19236
rect 9508 19196 10232 19224
rect 7892 19184 7898 19196
rect 10226 19184 10232 19196
rect 10284 19184 10290 19236
rect 1486 19116 1492 19168
rect 1544 19116 1550 19168
rect 5537 19159 5595 19165
rect 5537 19125 5549 19159
rect 5583 19156 5595 19159
rect 5902 19156 5908 19168
rect 5583 19128 5908 19156
rect 5583 19125 5595 19128
rect 5537 19119 5595 19125
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 7374 19116 7380 19168
rect 7432 19156 7438 19168
rect 7745 19159 7803 19165
rect 7745 19156 7757 19159
rect 7432 19128 7757 19156
rect 7432 19116 7438 19128
rect 7745 19125 7757 19128
rect 7791 19125 7803 19159
rect 7745 19119 7803 19125
rect 8386 19116 8392 19168
rect 8444 19116 8450 19168
rect 9766 19116 9772 19168
rect 9824 19116 9830 19168
rect 10962 19116 10968 19168
rect 11020 19116 11026 19168
rect 1104 19066 22356 19088
rect 1104 19014 3606 19066
rect 3658 19014 3670 19066
rect 3722 19014 3734 19066
rect 3786 19014 3798 19066
rect 3850 19014 3862 19066
rect 3914 19014 8919 19066
rect 8971 19014 8983 19066
rect 9035 19014 9047 19066
rect 9099 19014 9111 19066
rect 9163 19014 9175 19066
rect 9227 19014 14232 19066
rect 14284 19014 14296 19066
rect 14348 19014 14360 19066
rect 14412 19014 14424 19066
rect 14476 19014 14488 19066
rect 14540 19014 19545 19066
rect 19597 19014 19609 19066
rect 19661 19014 19673 19066
rect 19725 19014 19737 19066
rect 19789 19014 19801 19066
rect 19853 19014 22356 19066
rect 1104 18992 22356 19014
rect 4982 18912 4988 18964
rect 5040 18952 5046 18964
rect 5077 18955 5135 18961
rect 5077 18952 5089 18955
rect 5040 18924 5089 18952
rect 5040 18912 5046 18924
rect 5077 18921 5089 18924
rect 5123 18921 5135 18955
rect 5077 18915 5135 18921
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18952 6515 18955
rect 7834 18952 7840 18964
rect 6503 18924 7840 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 2498 18816 2504 18828
rect 2424 18788 2504 18816
rect 842 18708 848 18760
rect 900 18748 906 18760
rect 2424 18757 2452 18788
rect 2498 18776 2504 18788
rect 2556 18816 2562 18828
rect 2869 18819 2927 18825
rect 2869 18816 2881 18819
rect 2556 18788 2881 18816
rect 2556 18776 2562 18788
rect 2869 18785 2881 18788
rect 2915 18816 2927 18819
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 2915 18788 4261 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18816 6239 18819
rect 6472 18816 6500 18915
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 10045 18955 10103 18961
rect 10045 18921 10057 18955
rect 10091 18952 10103 18955
rect 10134 18952 10140 18964
rect 10091 18924 10140 18952
rect 10091 18921 10103 18924
rect 10045 18915 10103 18921
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 6638 18844 6644 18896
rect 6696 18884 6702 18896
rect 14090 18884 14096 18896
rect 6696 18856 14096 18884
rect 6696 18844 6702 18856
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 6227 18788 6500 18816
rect 6227 18785 6239 18788
rect 6181 18779 6239 18785
rect 8386 18776 8392 18828
rect 8444 18776 8450 18828
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 8628 18788 9904 18816
rect 8628 18776 8634 18788
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 900 18720 1409 18748
rect 900 18708 906 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18717 2467 18751
rect 2409 18711 2467 18717
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18748 2651 18751
rect 2958 18748 2964 18760
rect 2639 18720 2964 18748
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 2958 18708 2964 18720
rect 3016 18748 3022 18760
rect 3053 18751 3111 18757
rect 3053 18748 3065 18751
rect 3016 18720 3065 18748
rect 3016 18708 3022 18720
rect 3053 18717 3065 18720
rect 3099 18748 3111 18751
rect 4433 18751 4491 18757
rect 4433 18748 4445 18751
rect 3099 18720 4445 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 4433 18717 4445 18720
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 5166 18708 5172 18760
rect 5224 18708 5230 18760
rect 5902 18708 5908 18760
rect 5960 18708 5966 18760
rect 5997 18751 6055 18757
rect 5997 18717 6009 18751
rect 6043 18748 6055 18751
rect 6733 18751 6791 18757
rect 6733 18748 6745 18751
rect 6043 18720 6745 18748
rect 6043 18717 6055 18720
rect 5997 18711 6055 18717
rect 6733 18717 6745 18720
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 9766 18748 9772 18760
rect 8343 18720 9772 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 3237 18683 3295 18689
rect 3237 18649 3249 18683
rect 3283 18680 3295 18683
rect 4709 18683 4767 18689
rect 4709 18680 4721 18683
rect 3283 18652 4721 18680
rect 3283 18649 3295 18652
rect 3237 18643 3295 18649
rect 4709 18649 4721 18652
rect 4755 18649 4767 18683
rect 4709 18643 4767 18649
rect 4798 18640 4804 18692
rect 4856 18680 4862 18692
rect 4893 18683 4951 18689
rect 4893 18680 4905 18683
rect 4856 18652 4905 18680
rect 4856 18640 4862 18652
rect 4893 18649 4905 18652
rect 4939 18649 4951 18683
rect 4893 18643 4951 18649
rect 6546 18640 6552 18692
rect 6604 18640 6610 18692
rect 9876 18680 9904 18788
rect 10410 18776 10416 18828
rect 10468 18776 10474 18828
rect 10226 18708 10232 18760
rect 10284 18708 10290 18760
rect 18138 18708 18144 18760
rect 18196 18708 18202 18760
rect 22002 18708 22008 18760
rect 22060 18708 22066 18760
rect 12526 18680 12532 18692
rect 9876 18652 12532 18680
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 1854 18612 1860 18624
rect 1627 18584 1860 18612
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 1854 18572 1860 18584
rect 1912 18572 1918 18624
rect 2774 18572 2780 18624
rect 2832 18572 2838 18624
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 4617 18615 4675 18621
rect 4617 18612 4629 18615
rect 3384 18584 4629 18612
rect 3384 18572 3390 18584
rect 4617 18581 4629 18584
rect 4663 18581 4675 18615
rect 4617 18575 4675 18581
rect 5537 18615 5595 18621
rect 5537 18581 5549 18615
rect 5583 18612 5595 18615
rect 5626 18612 5632 18624
rect 5583 18584 5632 18612
rect 5583 18581 5595 18584
rect 5537 18575 5595 18581
rect 5626 18572 5632 18584
rect 5684 18572 5690 18624
rect 7558 18572 7564 18624
rect 7616 18612 7622 18624
rect 7929 18615 7987 18621
rect 7929 18612 7941 18615
rect 7616 18584 7941 18612
rect 7616 18572 7622 18584
rect 7929 18581 7941 18584
rect 7975 18581 7987 18615
rect 7929 18575 7987 18581
rect 20990 18572 20996 18624
rect 21048 18612 21054 18624
rect 21821 18615 21879 18621
rect 21821 18612 21833 18615
rect 21048 18584 21833 18612
rect 21048 18572 21054 18584
rect 21821 18581 21833 18584
rect 21867 18581 21879 18615
rect 21821 18575 21879 18581
rect 1104 18522 22356 18544
rect 1104 18470 4266 18522
rect 4318 18470 4330 18522
rect 4382 18470 4394 18522
rect 4446 18470 4458 18522
rect 4510 18470 4522 18522
rect 4574 18470 9579 18522
rect 9631 18470 9643 18522
rect 9695 18470 9707 18522
rect 9759 18470 9771 18522
rect 9823 18470 9835 18522
rect 9887 18470 14892 18522
rect 14944 18470 14956 18522
rect 15008 18470 15020 18522
rect 15072 18470 15084 18522
rect 15136 18470 15148 18522
rect 15200 18470 20205 18522
rect 20257 18470 20269 18522
rect 20321 18470 20333 18522
rect 20385 18470 20397 18522
rect 20449 18470 20461 18522
rect 20513 18470 22356 18522
rect 1104 18448 22356 18470
rect 1578 18368 1584 18420
rect 1636 18408 1642 18420
rect 2501 18411 2559 18417
rect 2501 18408 2513 18411
rect 1636 18380 2513 18408
rect 1636 18368 1642 18380
rect 2501 18377 2513 18380
rect 2547 18408 2559 18411
rect 2590 18408 2596 18420
rect 2547 18380 2596 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 3237 18411 3295 18417
rect 3237 18408 3249 18411
rect 2832 18380 3249 18408
rect 2832 18368 2838 18380
rect 3237 18377 3249 18380
rect 3283 18377 3295 18411
rect 3237 18371 3295 18377
rect 3326 18368 3332 18420
rect 3384 18368 3390 18420
rect 4264 18380 4936 18408
rect 4264 18340 4292 18380
rect 1688 18312 4292 18340
rect 4341 18343 4399 18349
rect 1688 18281 1716 18312
rect 4341 18309 4353 18343
rect 4387 18340 4399 18343
rect 4798 18340 4804 18352
rect 4387 18312 4804 18340
rect 4387 18309 4399 18312
rect 4341 18303 4399 18309
rect 4798 18300 4804 18312
rect 4856 18300 4862 18352
rect 4908 18340 4936 18380
rect 5626 18368 5632 18420
rect 5684 18368 5690 18420
rect 5718 18368 5724 18420
rect 5776 18368 5782 18420
rect 7190 18368 7196 18420
rect 7248 18368 7254 18420
rect 7745 18411 7803 18417
rect 7745 18377 7757 18411
rect 7791 18408 7803 18411
rect 7926 18408 7932 18420
rect 7791 18380 7932 18408
rect 7791 18377 7803 18380
rect 7745 18371 7803 18377
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 13538 18368 13544 18420
rect 13596 18368 13602 18420
rect 16025 18411 16083 18417
rect 16025 18377 16037 18411
rect 16071 18408 16083 18411
rect 16666 18408 16672 18420
rect 16071 18380 16672 18408
rect 16071 18377 16083 18380
rect 16025 18371 16083 18377
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 17313 18411 17371 18417
rect 17313 18377 17325 18411
rect 17359 18408 17371 18411
rect 17681 18411 17739 18417
rect 17681 18408 17693 18411
rect 17359 18380 17693 18408
rect 17359 18377 17371 18380
rect 17313 18371 17371 18377
rect 17681 18377 17693 18380
rect 17727 18377 17739 18411
rect 17681 18371 17739 18377
rect 18138 18368 18144 18420
rect 18196 18368 18202 18420
rect 18693 18411 18751 18417
rect 18693 18377 18705 18411
rect 18739 18377 18751 18411
rect 19981 18411 20039 18417
rect 19981 18408 19993 18411
rect 18693 18371 18751 18377
rect 19904 18380 19993 18408
rect 6914 18340 6920 18352
rect 4908 18312 6920 18340
rect 6914 18300 6920 18312
rect 6972 18300 6978 18352
rect 13814 18300 13820 18352
rect 13872 18340 13878 18352
rect 14001 18343 14059 18349
rect 14001 18340 14013 18343
rect 13872 18312 14013 18340
rect 13872 18300 13878 18312
rect 14001 18309 14013 18312
rect 14047 18309 14059 18343
rect 14001 18303 14059 18309
rect 14090 18300 14096 18352
rect 14148 18340 14154 18352
rect 17034 18340 17040 18352
rect 14148 18312 17040 18340
rect 14148 18300 14154 18312
rect 17034 18300 17040 18312
rect 17092 18300 17098 18352
rect 17221 18343 17279 18349
rect 17221 18309 17233 18343
rect 17267 18340 17279 18343
rect 18708 18340 18736 18371
rect 19904 18352 19932 18380
rect 19981 18377 19993 18380
rect 20027 18377 20039 18411
rect 19981 18371 20039 18377
rect 17267 18312 18736 18340
rect 19061 18343 19119 18349
rect 17267 18309 17279 18312
rect 17221 18303 17279 18309
rect 19061 18309 19073 18343
rect 19107 18340 19119 18343
rect 19334 18340 19340 18352
rect 19107 18312 19340 18340
rect 19107 18309 19119 18312
rect 19061 18303 19119 18309
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 19426 18300 19432 18352
rect 19484 18340 19490 18352
rect 19705 18343 19763 18349
rect 19705 18340 19717 18343
rect 19484 18312 19717 18340
rect 19484 18300 19490 18312
rect 19705 18309 19717 18312
rect 19751 18309 19763 18343
rect 19705 18303 19763 18309
rect 19886 18300 19892 18352
rect 19944 18300 19950 18352
rect 20349 18343 20407 18349
rect 20349 18309 20361 18343
rect 20395 18340 20407 18343
rect 20395 18312 21036 18340
rect 20395 18309 20407 18312
rect 20349 18303 20407 18309
rect 21008 18284 21036 18312
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 1854 18232 1860 18284
rect 1912 18281 1918 18284
rect 1912 18275 1950 18281
rect 1938 18241 1950 18275
rect 2866 18272 2872 18284
rect 1912 18235 1950 18241
rect 2746 18244 2872 18272
rect 1912 18232 1918 18235
rect 2317 18207 2375 18213
rect 2317 18173 2329 18207
rect 2363 18173 2375 18207
rect 2317 18167 2375 18173
rect 2332 18136 2360 18167
rect 2406 18164 2412 18216
rect 2464 18164 2470 18216
rect 2746 18136 2774 18244
rect 2866 18232 2872 18244
rect 2924 18232 2930 18284
rect 3881 18275 3939 18281
rect 3881 18241 3893 18275
rect 3927 18272 3939 18275
rect 4062 18272 4068 18284
rect 3927 18244 4068 18272
rect 3927 18241 3939 18244
rect 3881 18235 3939 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4890 18232 4896 18284
rect 4948 18272 4954 18284
rect 5718 18272 5724 18284
rect 4948 18244 5724 18272
rect 4948 18232 4954 18244
rect 5718 18232 5724 18244
rect 5776 18272 5782 18284
rect 6638 18272 6644 18284
rect 5776 18244 6644 18272
rect 5776 18232 5782 18244
rect 6638 18232 6644 18244
rect 6696 18232 6702 18284
rect 7374 18232 7380 18284
rect 7432 18232 7438 18284
rect 7558 18232 7564 18284
rect 7616 18232 7622 18284
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 13173 18275 13231 18281
rect 13173 18272 13185 18275
rect 13127 18244 13185 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 13173 18241 13185 18244
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 13354 18232 13360 18284
rect 13412 18232 13418 18284
rect 13630 18232 13636 18284
rect 13688 18232 13694 18284
rect 13906 18232 13912 18284
rect 13964 18232 13970 18284
rect 15838 18232 15844 18284
rect 15896 18232 15902 18284
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18241 16175 18275
rect 16117 18235 16175 18241
rect 3145 18207 3203 18213
rect 3145 18173 3157 18207
rect 3191 18173 3203 18207
rect 3145 18167 3203 18173
rect 3789 18207 3847 18213
rect 3789 18173 3801 18207
rect 3835 18204 3847 18207
rect 3970 18204 3976 18216
rect 3835 18176 3976 18204
rect 3835 18173 3847 18176
rect 3789 18167 3847 18173
rect 2332 18108 2774 18136
rect 2869 18139 2927 18145
rect 2869 18105 2881 18139
rect 2915 18136 2927 18139
rect 2958 18136 2964 18148
rect 2915 18108 2964 18136
rect 2915 18105 2927 18108
rect 2869 18099 2927 18105
rect 2958 18096 2964 18108
rect 3016 18096 3022 18148
rect 1486 18028 1492 18080
rect 1544 18028 1550 18080
rect 1946 18028 1952 18080
rect 2004 18077 2010 18080
rect 2004 18071 2053 18077
rect 2004 18037 2007 18071
rect 2041 18037 2053 18071
rect 3160 18068 3188 18167
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 5169 18207 5227 18213
rect 5169 18173 5181 18207
rect 5215 18204 5227 18207
rect 5537 18207 5595 18213
rect 5537 18204 5549 18207
rect 5215 18176 5549 18204
rect 5215 18173 5227 18176
rect 5169 18167 5227 18173
rect 5537 18173 5549 18176
rect 5583 18204 5595 18207
rect 5810 18204 5816 18216
rect 5583 18176 5816 18204
rect 5583 18173 5595 18176
rect 5537 18167 5595 18173
rect 5810 18164 5816 18176
rect 5868 18164 5874 18216
rect 12894 18164 12900 18216
rect 12952 18164 12958 18216
rect 3697 18139 3755 18145
rect 3697 18105 3709 18139
rect 3743 18136 3755 18139
rect 5994 18136 6000 18148
rect 3743 18108 6000 18136
rect 3743 18105 3755 18108
rect 3697 18099 3755 18105
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 12710 18096 12716 18148
rect 12768 18096 12774 18148
rect 13262 18096 13268 18148
rect 13320 18136 13326 18148
rect 13633 18139 13691 18145
rect 13633 18136 13645 18139
rect 13320 18108 13645 18136
rect 13320 18096 13326 18108
rect 13633 18105 13645 18108
rect 13679 18105 13691 18139
rect 13633 18099 13691 18105
rect 13817 18139 13875 18145
rect 13817 18105 13829 18139
rect 13863 18136 13875 18139
rect 16132 18136 16160 18235
rect 18046 18232 18052 18284
rect 18104 18232 18110 18284
rect 20990 18281 20996 18284
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18272 19211 18275
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19199 18244 19533 18272
rect 19199 18241 19211 18244
rect 19153 18235 19211 18241
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18272 20499 18275
rect 20855 18275 20913 18281
rect 20855 18272 20867 18275
rect 20487 18244 20867 18272
rect 20487 18241 20499 18244
rect 20441 18235 20499 18241
rect 20855 18241 20867 18244
rect 20901 18241 20913 18275
rect 20855 18235 20913 18241
rect 20958 18275 20996 18281
rect 20958 18241 20970 18275
rect 20958 18235 20996 18241
rect 20990 18232 20996 18235
rect 21048 18232 21054 18284
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 21361 18275 21419 18281
rect 21361 18272 21373 18275
rect 21140 18244 21373 18272
rect 21140 18232 21146 18244
rect 21361 18241 21373 18244
rect 21407 18241 21419 18275
rect 21361 18235 21419 18241
rect 17402 18164 17408 18216
rect 17460 18164 17466 18216
rect 18325 18207 18383 18213
rect 18325 18173 18337 18207
rect 18371 18204 18383 18207
rect 18414 18204 18420 18216
rect 18371 18176 18420 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 18414 18164 18420 18176
rect 18472 18204 18478 18216
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 18472 18176 19257 18204
rect 18472 18164 18478 18176
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19245 18167 19303 18173
rect 20530 18164 20536 18216
rect 20588 18164 20594 18216
rect 13863 18108 16160 18136
rect 13863 18105 13875 18108
rect 13817 18099 13875 18105
rect 4154 18068 4160 18080
rect 3160 18040 4160 18068
rect 2004 18031 2053 18037
rect 2004 18028 2010 18031
rect 4154 18028 4160 18040
rect 4212 18068 4218 18080
rect 4890 18068 4896 18080
rect 4212 18040 4896 18068
rect 4212 18028 4218 18040
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 6089 18071 6147 18077
rect 6089 18037 6101 18071
rect 6135 18068 6147 18071
rect 6178 18068 6184 18080
rect 6135 18040 6184 18068
rect 6135 18037 6147 18040
rect 6089 18031 6147 18037
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 16132 18068 16160 18108
rect 16301 18139 16359 18145
rect 16301 18105 16313 18139
rect 16347 18136 16359 18139
rect 17310 18136 17316 18148
rect 16347 18108 17316 18136
rect 16347 18105 16359 18108
rect 16301 18099 16359 18105
rect 17310 18096 17316 18108
rect 17368 18096 17374 18148
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 16132 18040 16865 18068
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 21542 18028 21548 18080
rect 21600 18028 21606 18080
rect 1104 17978 22356 18000
rect 1104 17926 3606 17978
rect 3658 17926 3670 17978
rect 3722 17926 3734 17978
rect 3786 17926 3798 17978
rect 3850 17926 3862 17978
rect 3914 17926 8919 17978
rect 8971 17926 8983 17978
rect 9035 17926 9047 17978
rect 9099 17926 9111 17978
rect 9163 17926 9175 17978
rect 9227 17926 14232 17978
rect 14284 17926 14296 17978
rect 14348 17926 14360 17978
rect 14412 17926 14424 17978
rect 14476 17926 14488 17978
rect 14540 17926 19545 17978
rect 19597 17926 19609 17978
rect 19661 17926 19673 17978
rect 19725 17926 19737 17978
rect 19789 17926 19801 17978
rect 19853 17926 22356 17978
rect 1104 17904 22356 17926
rect 2406 17824 2412 17876
rect 2464 17864 2470 17876
rect 2547 17867 2605 17873
rect 2547 17864 2559 17867
rect 2464 17836 2559 17864
rect 2464 17824 2470 17836
rect 2547 17833 2559 17836
rect 2593 17833 2605 17867
rect 4706 17864 4712 17876
rect 2547 17827 2605 17833
rect 2884 17836 4712 17864
rect 2884 17796 2912 17836
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 6914 17824 6920 17876
rect 6972 17824 6978 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7469 17867 7527 17873
rect 7469 17864 7481 17867
rect 7432 17836 7481 17864
rect 7432 17824 7438 17836
rect 7469 17833 7481 17836
rect 7515 17833 7527 17867
rect 7469 17827 7527 17833
rect 12253 17867 12311 17873
rect 12253 17833 12265 17867
rect 12299 17864 12311 17867
rect 13354 17864 13360 17876
rect 12299 17836 13360 17864
rect 12299 17833 12311 17836
rect 12253 17827 12311 17833
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 18046 17824 18052 17876
rect 18104 17824 18110 17876
rect 1780 17768 2912 17796
rect 1780 17740 1808 17768
rect 2958 17756 2964 17808
rect 3016 17796 3022 17808
rect 3016 17768 3096 17796
rect 3016 17756 3022 17768
rect 1762 17688 1768 17740
rect 1820 17688 1826 17740
rect 1946 17688 1952 17740
rect 2004 17688 2010 17740
rect 3068 17737 3096 17768
rect 4062 17756 4068 17808
rect 4120 17756 4126 17808
rect 13173 17799 13231 17805
rect 13173 17796 13185 17799
rect 12452 17768 13185 17796
rect 3053 17731 3111 17737
rect 3053 17697 3065 17731
rect 3099 17697 3111 17731
rect 3053 17691 3111 17697
rect 3329 17731 3387 17737
rect 3329 17697 3341 17731
rect 3375 17728 3387 17731
rect 4080 17728 4108 17756
rect 4157 17731 4215 17737
rect 4157 17728 4169 17731
rect 3375 17700 4169 17728
rect 3375 17697 3387 17700
rect 3329 17691 3387 17697
rect 4157 17697 4169 17700
rect 4203 17697 4215 17731
rect 4157 17691 4215 17697
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 1854 17620 1860 17672
rect 1912 17660 1918 17672
rect 2041 17663 2099 17669
rect 2041 17660 2053 17663
rect 1912 17632 2053 17660
rect 1912 17620 1918 17632
rect 2041 17629 2053 17632
rect 2087 17629 2099 17663
rect 2041 17623 2099 17629
rect 2590 17620 2596 17672
rect 2648 17669 2654 17672
rect 2648 17663 2676 17669
rect 2664 17629 2676 17663
rect 2648 17623 2676 17629
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 2648 17620 2654 17623
rect 2976 17592 3004 17623
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 4028 17632 4077 17660
rect 4028 17620 4034 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 2746 17564 3004 17592
rect 4448 17592 4476 17691
rect 4890 17688 4896 17740
rect 4948 17688 4954 17740
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17728 5135 17731
rect 5166 17728 5172 17740
rect 5123 17700 5172 17728
rect 5123 17697 5135 17700
rect 5077 17691 5135 17697
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 5810 17688 5816 17740
rect 5868 17688 5874 17740
rect 8846 17688 8852 17740
rect 8904 17728 8910 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 8904 17700 9873 17728
rect 8904 17688 8910 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 10134 17688 10140 17740
rect 10192 17688 10198 17740
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17728 10563 17731
rect 10962 17728 10968 17740
rect 10551 17700 10968 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 5994 17620 6000 17672
rect 6052 17620 6058 17672
rect 7101 17663 7159 17669
rect 7101 17660 7113 17663
rect 6886 17632 7113 17660
rect 5169 17595 5227 17601
rect 5169 17592 5181 17595
rect 4448 17564 5181 17592
rect 2409 17527 2467 17533
rect 2409 17493 2421 17527
rect 2455 17524 2467 17527
rect 2498 17524 2504 17536
rect 2455 17496 2504 17524
rect 2455 17493 2467 17496
rect 2409 17487 2467 17493
rect 2498 17484 2504 17496
rect 2556 17524 2562 17536
rect 2746 17524 2774 17564
rect 5169 17561 5181 17564
rect 5215 17561 5227 17595
rect 5169 17555 5227 17561
rect 2556 17496 2774 17524
rect 5537 17527 5595 17533
rect 2556 17484 2562 17496
rect 5537 17493 5549 17527
rect 5583 17524 5595 17527
rect 5905 17527 5963 17533
rect 5905 17524 5917 17527
rect 5583 17496 5917 17524
rect 5583 17493 5595 17496
rect 5537 17487 5595 17493
rect 5905 17493 5917 17496
rect 5951 17493 5963 17527
rect 5905 17487 5963 17493
rect 6365 17527 6423 17533
rect 6365 17493 6377 17527
rect 6411 17524 6423 17527
rect 6886 17524 6914 17632
rect 7101 17629 7113 17632
rect 7147 17660 7159 17663
rect 7377 17663 7435 17669
rect 7377 17660 7389 17663
rect 7147 17632 7389 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 7377 17629 7389 17632
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 7653 17663 7711 17669
rect 7653 17660 7665 17663
rect 7616 17632 7665 17660
rect 7616 17620 7622 17632
rect 7653 17629 7665 17632
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 8938 17620 8944 17672
rect 8996 17620 9002 17672
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17660 10287 17663
rect 10520 17660 10548 17691
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 12452 17669 12480 17768
rect 13173 17765 13185 17768
rect 13219 17796 13231 17799
rect 13219 17768 13400 17796
rect 13219 17765 13231 17768
rect 13173 17759 13231 17765
rect 12529 17731 12587 17737
rect 12529 17697 12541 17731
rect 12575 17697 12587 17731
rect 12529 17691 12587 17697
rect 10275 17632 10548 17660
rect 10597 17663 10655 17669
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 10597 17629 10609 17663
rect 10643 17629 10655 17663
rect 10597 17623 10655 17629
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17660 11115 17663
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 11103 17632 11345 17660
rect 11103 17629 11115 17632
rect 11057 17623 11115 17629
rect 11333 17629 11345 17632
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 7285 17595 7343 17601
rect 7285 17561 7297 17595
rect 7331 17592 7343 17595
rect 7742 17592 7748 17604
rect 7331 17564 7748 17592
rect 7331 17561 7343 17564
rect 7285 17555 7343 17561
rect 7742 17552 7748 17564
rect 7800 17552 7806 17604
rect 10134 17552 10140 17604
rect 10192 17592 10198 17604
rect 10612 17592 10640 17623
rect 10192 17564 10640 17592
rect 10192 17552 10198 17564
rect 11146 17552 11152 17604
rect 11204 17552 11210 17604
rect 11517 17595 11575 17601
rect 11517 17561 11529 17595
rect 11563 17592 11575 17595
rect 12544 17592 12572 17691
rect 12894 17688 12900 17740
rect 12952 17688 12958 17740
rect 13372 17737 13400 17768
rect 13446 17756 13452 17808
rect 13504 17796 13510 17808
rect 20165 17799 20223 17805
rect 13504 17768 15608 17796
rect 13504 17756 13510 17768
rect 15580 17737 15608 17768
rect 20165 17765 20177 17799
rect 20211 17765 20223 17799
rect 20165 17759 20223 17765
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 13817 17731 13875 17737
rect 13817 17697 13829 17731
rect 13863 17728 13875 17731
rect 15565 17731 15623 17737
rect 13863 17700 15424 17728
rect 13863 17697 13875 17700
rect 13817 17691 13875 17697
rect 12710 17620 12716 17672
rect 12768 17660 12774 17672
rect 15396 17669 15424 17700
rect 15565 17697 15577 17731
rect 15611 17728 15623 17731
rect 16390 17728 16396 17740
rect 15611 17700 16396 17728
rect 15611 17697 15623 17700
rect 15565 17691 15623 17697
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 18325 17731 18383 17737
rect 18325 17697 18337 17731
rect 18371 17728 18383 17731
rect 18598 17728 18604 17740
rect 18371 17700 18604 17728
rect 18371 17697 18383 17700
rect 18325 17691 18383 17697
rect 18598 17688 18604 17700
rect 18656 17728 18662 17740
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 18656 17700 19257 17728
rect 18656 17688 18662 17700
rect 19245 17697 19257 17700
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 19518 17688 19524 17740
rect 19576 17728 19582 17740
rect 20180 17728 20208 17759
rect 19576 17700 20208 17728
rect 19576 17688 19582 17700
rect 20622 17688 20628 17740
rect 20680 17728 20686 17740
rect 20717 17731 20775 17737
rect 20717 17728 20729 17731
rect 20680 17700 20729 17728
rect 20680 17688 20686 17700
rect 20717 17697 20729 17700
rect 20763 17697 20775 17731
rect 20717 17691 20775 17697
rect 12805 17663 12863 17669
rect 12805 17660 12817 17663
rect 12768 17632 12817 17660
rect 12768 17620 12774 17632
rect 12805 17629 12817 17632
rect 12851 17629 12863 17663
rect 12805 17623 12863 17629
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17629 15439 17663
rect 15381 17623 15439 17629
rect 15473 17663 15531 17669
rect 15473 17629 15485 17663
rect 15519 17660 15531 17663
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15519 17632 15853 17660
rect 15519 17629 15531 17632
rect 15473 17623 15531 17629
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 18506 17660 18512 17672
rect 18463 17632 18512 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 13464 17592 13492 17623
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19886 17660 19892 17672
rect 19659 17632 19892 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17660 20591 17663
rect 21142 17663 21200 17669
rect 21142 17660 21154 17663
rect 20579 17632 21154 17660
rect 20579 17629 20591 17632
rect 20533 17623 20591 17629
rect 21142 17629 21154 17632
rect 21188 17660 21200 17663
rect 21818 17660 21824 17672
rect 21188 17632 21824 17660
rect 21188 17629 21200 17632
rect 21142 17623 21200 17629
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 11563 17564 13492 17592
rect 11563 17561 11575 17564
rect 11517 17555 11575 17561
rect 18782 17552 18788 17604
rect 18840 17592 18846 17604
rect 18877 17595 18935 17601
rect 18877 17592 18889 17595
rect 18840 17564 18889 17592
rect 18840 17552 18846 17564
rect 18877 17561 18889 17564
rect 18923 17561 18935 17595
rect 18877 17555 18935 17561
rect 19058 17552 19064 17604
rect 19116 17552 19122 17604
rect 6411 17496 6914 17524
rect 7561 17527 7619 17533
rect 6411 17493 6423 17496
rect 6365 17487 6423 17493
rect 7561 17493 7573 17527
rect 7607 17524 7619 17527
rect 8662 17524 8668 17536
rect 7607 17496 8668 17524
rect 7607 17493 7619 17496
rect 7561 17487 7619 17493
rect 8662 17484 8668 17496
rect 8720 17484 8726 17536
rect 15013 17527 15071 17533
rect 15013 17493 15025 17527
rect 15059 17524 15071 17527
rect 15286 17524 15292 17536
rect 15059 17496 15292 17524
rect 15059 17493 15071 17496
rect 15013 17487 15071 17493
rect 15286 17484 15292 17496
rect 15344 17484 15350 17536
rect 18690 17484 18696 17536
rect 18748 17484 18754 17536
rect 20625 17527 20683 17533
rect 20625 17493 20637 17527
rect 20671 17524 20683 17527
rect 21039 17527 21097 17533
rect 21039 17524 21051 17527
rect 20671 17496 21051 17524
rect 20671 17493 20683 17496
rect 20625 17487 20683 17493
rect 21039 17493 21051 17496
rect 21085 17493 21097 17527
rect 21039 17487 21097 17493
rect 1104 17434 22356 17456
rect 1104 17382 4266 17434
rect 4318 17382 4330 17434
rect 4382 17382 4394 17434
rect 4446 17382 4458 17434
rect 4510 17382 4522 17434
rect 4574 17382 9579 17434
rect 9631 17382 9643 17434
rect 9695 17382 9707 17434
rect 9759 17382 9771 17434
rect 9823 17382 9835 17434
rect 9887 17382 14892 17434
rect 14944 17382 14956 17434
rect 15008 17382 15020 17434
rect 15072 17382 15084 17434
rect 15136 17382 15148 17434
rect 15200 17382 20205 17434
rect 20257 17382 20269 17434
rect 20321 17382 20333 17434
rect 20385 17382 20397 17434
rect 20449 17382 20461 17434
rect 20513 17382 22356 17434
rect 1104 17360 22356 17382
rect 5997 17323 6055 17329
rect 5997 17289 6009 17323
rect 6043 17289 6055 17323
rect 5997 17283 6055 17289
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 6012 17184 6040 17283
rect 8846 17280 8852 17332
rect 8904 17280 8910 17332
rect 8938 17280 8944 17332
rect 8996 17280 9002 17332
rect 11057 17323 11115 17329
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 11146 17320 11152 17332
rect 11103 17292 11152 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 14277 17323 14335 17329
rect 14277 17289 14289 17323
rect 14323 17289 14335 17323
rect 14277 17283 14335 17289
rect 15105 17323 15163 17329
rect 15105 17289 15117 17323
rect 15151 17320 15163 17323
rect 15286 17320 15292 17332
rect 15151 17292 15292 17320
rect 15151 17289 15163 17292
rect 15105 17283 15163 17289
rect 10502 17212 10508 17264
rect 10560 17252 10566 17264
rect 12621 17255 12679 17261
rect 10560 17224 10916 17252
rect 10560 17212 10566 17224
rect 1719 17156 6040 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 6178 17144 6184 17196
rect 6236 17144 6242 17196
rect 10888 17193 10916 17224
rect 12621 17221 12633 17255
rect 12667 17252 12679 17255
rect 12710 17252 12716 17264
rect 12667 17224 12716 17252
rect 12667 17221 12679 17224
rect 12621 17215 12679 17221
rect 12710 17212 12716 17224
rect 12768 17212 12774 17264
rect 12805 17255 12863 17261
rect 12805 17221 12817 17255
rect 12851 17252 12863 17255
rect 12894 17252 12900 17264
rect 12851 17224 12900 17252
rect 12851 17221 12863 17224
rect 12805 17215 12863 17221
rect 12894 17212 12900 17224
rect 12952 17212 12958 17264
rect 12989 17255 13047 17261
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 13817 17255 13875 17261
rect 13817 17252 13829 17255
rect 13035 17224 13829 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 13817 17221 13829 17224
rect 13863 17221 13875 17255
rect 14292 17252 14320 17283
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 15565 17323 15623 17329
rect 15565 17289 15577 17323
rect 15611 17289 15623 17323
rect 15565 17283 15623 17289
rect 15841 17323 15899 17329
rect 15841 17289 15853 17323
rect 15887 17320 15899 17323
rect 17954 17320 17960 17332
rect 15887 17292 17960 17320
rect 15887 17289 15899 17292
rect 15841 17283 15899 17289
rect 15197 17255 15255 17261
rect 15197 17252 15209 17255
rect 14292 17224 15209 17252
rect 13817 17215 13875 17221
rect 15197 17221 15209 17224
rect 15243 17221 15255 17255
rect 15197 17215 15255 17221
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 10873 17187 10931 17193
rect 10459 17156 10732 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 9033 17119 9091 17125
rect 9033 17116 9045 17119
rect 8536 17088 9045 17116
rect 8536 17076 8542 17088
rect 9033 17085 9045 17088
rect 9079 17085 9091 17119
rect 9033 17079 9091 17085
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 10134 17116 10140 17128
rect 10091 17088 10140 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 10502 17076 10508 17128
rect 10560 17076 10566 17128
rect 842 17008 848 17060
rect 900 17048 906 17060
rect 10704 17057 10732 17156
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 12728 17116 12756 17212
rect 12912 17184 12940 17212
rect 13265 17187 13323 17193
rect 13265 17184 13277 17187
rect 12912 17156 13277 17184
rect 13265 17153 13277 17156
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17184 13507 17187
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 13495 17156 13921 17184
rect 13495 17153 13507 17156
rect 13449 17147 13507 17153
rect 13909 17153 13921 17156
rect 13955 17153 13967 17187
rect 15580 17184 15608 17283
rect 17954 17280 17960 17292
rect 18012 17280 18018 17332
rect 18782 17280 18788 17332
rect 18840 17280 18846 17332
rect 18877 17323 18935 17329
rect 18877 17289 18889 17323
rect 18923 17320 18935 17323
rect 19058 17320 19064 17332
rect 18923 17292 19064 17320
rect 18923 17289 18935 17292
rect 18877 17283 18935 17289
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19334 17280 19340 17332
rect 19392 17280 19398 17332
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 15580 17156 15669 17184
rect 13909 17147 13967 17153
rect 15657 17153 15669 17156
rect 15703 17184 15715 17187
rect 15746 17184 15752 17196
rect 15703 17156 15752 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 18598 17144 18604 17196
rect 18656 17144 18662 17196
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19518 17184 19524 17196
rect 19107 17156 19524 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 21358 17144 21364 17196
rect 21416 17144 21422 17196
rect 12986 17116 12992 17128
rect 12728 17088 12992 17116
rect 12986 17076 12992 17088
rect 13044 17116 13050 17128
rect 13081 17119 13139 17125
rect 13081 17116 13093 17119
rect 13044 17088 13093 17116
rect 13044 17076 13050 17088
rect 13081 17085 13093 17088
rect 13127 17085 13139 17119
rect 13081 17079 13139 17085
rect 13538 17076 13544 17128
rect 13596 17116 13602 17128
rect 13633 17119 13691 17125
rect 13633 17116 13645 17119
rect 13596 17088 13645 17116
rect 13596 17076 13602 17088
rect 13633 17085 13645 17088
rect 13679 17116 13691 17119
rect 13722 17116 13728 17128
rect 13679 17088 13728 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17116 18475 17119
rect 18506 17116 18512 17128
rect 18463 17088 18512 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 1489 17051 1547 17057
rect 1489 17048 1501 17051
rect 900 17020 1501 17048
rect 900 17008 906 17020
rect 1489 17017 1501 17020
rect 1535 17017 1547 17051
rect 1489 17011 1547 17017
rect 10689 17051 10747 17057
rect 10689 17017 10701 17051
rect 10735 17048 10747 17051
rect 10778 17048 10784 17060
rect 10735 17020 10784 17048
rect 10735 17017 10747 17020
rect 10689 17011 10747 17017
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 14936 17048 14964 17079
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 19886 17116 19892 17128
rect 19751 17088 19892 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 12584 17020 14964 17048
rect 19245 17051 19303 17057
rect 12584 17008 12590 17020
rect 19245 17017 19257 17051
rect 19291 17048 19303 17051
rect 19720 17048 19748 17079
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 19291 17020 19748 17048
rect 19291 17017 19303 17020
rect 19245 17011 19303 17017
rect 21542 17008 21548 17060
rect 21600 17008 21606 17060
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 8352 16952 8493 16980
rect 8352 16940 8358 16952
rect 8481 16949 8493 16952
rect 8527 16949 8539 16983
rect 8481 16943 8539 16949
rect 1104 16890 22356 16912
rect 1104 16838 3606 16890
rect 3658 16838 3670 16890
rect 3722 16838 3734 16890
rect 3786 16838 3798 16890
rect 3850 16838 3862 16890
rect 3914 16838 8919 16890
rect 8971 16838 8983 16890
rect 9035 16838 9047 16890
rect 9099 16838 9111 16890
rect 9163 16838 9175 16890
rect 9227 16838 14232 16890
rect 14284 16838 14296 16890
rect 14348 16838 14360 16890
rect 14412 16838 14424 16890
rect 14476 16838 14488 16890
rect 14540 16838 19545 16890
rect 19597 16838 19609 16890
rect 19661 16838 19673 16890
rect 19725 16838 19737 16890
rect 19789 16838 19801 16890
rect 19853 16838 22356 16890
rect 1104 16816 22356 16838
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 10744 16748 12480 16776
rect 10744 16736 10750 16748
rect 8478 16668 8484 16720
rect 8536 16708 8542 16720
rect 11149 16711 11207 16717
rect 11149 16708 11161 16711
rect 8536 16680 9674 16708
rect 8536 16668 8542 16680
rect 8294 16600 8300 16652
rect 8352 16600 8358 16652
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 8570 16640 8576 16652
rect 8435 16612 8576 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 8570 16600 8576 16612
rect 8628 16600 8634 16652
rect 842 16532 848 16584
rect 900 16572 906 16584
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 900 16544 1409 16572
rect 900 16532 906 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 5626 16532 5632 16584
rect 5684 16532 5690 16584
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16541 7251 16575
rect 7193 16535 7251 16541
rect 6730 16464 6736 16516
rect 6788 16504 6794 16516
rect 7208 16504 7236 16535
rect 7742 16532 7748 16584
rect 7800 16532 7806 16584
rect 9646 16581 9674 16680
rect 9968 16680 11161 16708
rect 9968 16649 9996 16680
rect 11149 16677 11161 16680
rect 11195 16677 11207 16711
rect 11149 16671 11207 16677
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 10502 16600 10508 16652
rect 10560 16600 10566 16652
rect 12452 16649 12480 16748
rect 12986 16736 12992 16788
rect 13044 16736 13050 16788
rect 15657 16779 15715 16785
rect 15657 16745 15669 16779
rect 15703 16776 15715 16779
rect 15838 16776 15844 16788
rect 15703 16748 15844 16776
rect 15703 16745 15715 16748
rect 15657 16739 15715 16745
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 12894 16668 12900 16720
rect 12952 16708 12958 16720
rect 13081 16711 13139 16717
rect 13081 16708 13093 16711
rect 12952 16680 13093 16708
rect 12952 16668 12958 16680
rect 13081 16677 13093 16680
rect 13127 16677 13139 16711
rect 13081 16671 13139 16677
rect 15565 16711 15623 16717
rect 15565 16677 15577 16711
rect 15611 16708 15623 16711
rect 16485 16711 16543 16717
rect 15611 16680 16344 16708
rect 15611 16677 15623 16680
rect 15565 16671 15623 16677
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 12437 16643 12495 16649
rect 10735 16612 10824 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 9646 16575 9706 16581
rect 9646 16544 9660 16575
rect 9648 16541 9660 16544
rect 9694 16541 9706 16575
rect 9648 16535 9706 16541
rect 10796 16516 10824 16612
rect 12437 16609 12449 16643
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 13170 16640 13176 16652
rect 12676 16612 13176 16640
rect 12676 16600 12682 16612
rect 13170 16600 13176 16612
rect 13228 16640 13234 16652
rect 13633 16643 13691 16649
rect 13633 16640 13645 16643
rect 13228 16612 13645 16640
rect 13228 16600 13234 16612
rect 13633 16609 13645 16612
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 15746 16600 15752 16652
rect 15804 16600 15810 16652
rect 16316 16584 16344 16680
rect 16485 16677 16497 16711
rect 16531 16677 16543 16711
rect 16485 16671 16543 16677
rect 13446 16532 13452 16584
rect 13504 16572 13510 16584
rect 15286 16572 15292 16584
rect 13504 16544 15292 16572
rect 13504 16532 13510 16544
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15396 16544 15853 16572
rect 15396 16516 15424 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 16298 16572 16304 16584
rect 16259 16544 16304 16572
rect 15841 16535 15899 16541
rect 16298 16532 16304 16544
rect 16356 16532 16362 16584
rect 16500 16572 16528 16671
rect 21082 16572 21088 16584
rect 16500 16544 21088 16572
rect 21082 16532 21088 16544
rect 21140 16532 21146 16584
rect 22002 16532 22008 16584
rect 22060 16532 22066 16584
rect 6788 16476 7880 16504
rect 6788 16464 6794 16476
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16436 1639 16439
rect 2038 16436 2044 16448
rect 1627 16408 2044 16436
rect 1627 16405 1639 16408
rect 1581 16399 1639 16405
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 7006 16396 7012 16448
rect 7064 16396 7070 16448
rect 7466 16396 7472 16448
rect 7524 16436 7530 16448
rect 7852 16445 7880 16476
rect 10778 16464 10784 16516
rect 10836 16464 10842 16516
rect 10965 16507 11023 16513
rect 10965 16473 10977 16507
rect 11011 16473 11023 16507
rect 10965 16467 11023 16473
rect 12621 16507 12679 16513
rect 12621 16473 12633 16507
rect 12667 16504 12679 16507
rect 13814 16504 13820 16516
rect 12667 16476 13820 16504
rect 12667 16473 12679 16476
rect 12621 16467 12679 16473
rect 7561 16439 7619 16445
rect 7561 16436 7573 16439
rect 7524 16408 7573 16436
rect 7524 16396 7530 16408
rect 7561 16405 7573 16408
rect 7607 16405 7619 16439
rect 7561 16399 7619 16405
rect 7837 16439 7895 16445
rect 7837 16405 7849 16439
rect 7883 16405 7895 16439
rect 7837 16399 7895 16405
rect 8205 16439 8263 16445
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 9493 16439 9551 16445
rect 9493 16436 9505 16439
rect 8251 16408 9505 16436
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 9493 16405 9505 16408
rect 9539 16405 9551 16439
rect 9493 16399 9551 16405
rect 9861 16439 9919 16445
rect 9861 16405 9873 16439
rect 9907 16436 9919 16439
rect 10321 16439 10379 16445
rect 10321 16436 10333 16439
rect 9907 16408 10333 16436
rect 9907 16405 9919 16408
rect 9861 16399 9919 16405
rect 10321 16405 10333 16408
rect 10367 16405 10379 16439
rect 10321 16399 10379 16405
rect 10502 16396 10508 16448
rect 10560 16436 10566 16448
rect 10980 16436 11008 16467
rect 13814 16464 13820 16476
rect 13872 16464 13878 16516
rect 15378 16464 15384 16516
rect 15436 16464 15442 16516
rect 21358 16504 21364 16516
rect 16040 16476 21364 16504
rect 10560 16408 11008 16436
rect 10560 16396 10566 16408
rect 12526 16396 12532 16448
rect 12584 16396 12590 16448
rect 13538 16396 13544 16448
rect 13596 16396 13602 16448
rect 15473 16439 15531 16445
rect 15473 16405 15485 16439
rect 15519 16436 15531 16439
rect 15562 16436 15568 16448
rect 15519 16408 15568 16436
rect 15519 16405 15531 16408
rect 15473 16399 15531 16405
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 16040 16445 16068 16476
rect 21358 16464 21364 16476
rect 21416 16464 21422 16516
rect 16025 16439 16083 16445
rect 16025 16405 16037 16439
rect 16071 16405 16083 16439
rect 16025 16399 16083 16405
rect 21726 16396 21732 16448
rect 21784 16436 21790 16448
rect 21821 16439 21879 16445
rect 21821 16436 21833 16439
rect 21784 16408 21833 16436
rect 21784 16396 21790 16408
rect 21821 16405 21833 16408
rect 21867 16405 21879 16439
rect 21821 16399 21879 16405
rect 1104 16346 22356 16368
rect 1104 16294 4266 16346
rect 4318 16294 4330 16346
rect 4382 16294 4394 16346
rect 4446 16294 4458 16346
rect 4510 16294 4522 16346
rect 4574 16294 9579 16346
rect 9631 16294 9643 16346
rect 9695 16294 9707 16346
rect 9759 16294 9771 16346
rect 9823 16294 9835 16346
rect 9887 16294 14892 16346
rect 14944 16294 14956 16346
rect 15008 16294 15020 16346
rect 15072 16294 15084 16346
rect 15136 16294 15148 16346
rect 15200 16294 20205 16346
rect 20257 16294 20269 16346
rect 20321 16294 20333 16346
rect 20385 16294 20397 16346
rect 20449 16294 20461 16346
rect 20513 16294 22356 16346
rect 1104 16272 22356 16294
rect 3970 16192 3976 16244
rect 4028 16192 4034 16244
rect 5626 16192 5632 16244
rect 5684 16232 5690 16244
rect 5721 16235 5779 16241
rect 5721 16232 5733 16235
rect 5684 16204 5733 16232
rect 5684 16192 5690 16204
rect 5721 16201 5733 16204
rect 5767 16201 5779 16235
rect 5721 16195 5779 16201
rect 6822 16192 6828 16244
rect 6880 16192 6886 16244
rect 10502 16192 10508 16244
rect 10560 16232 10566 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 10560 16204 10609 16232
rect 10560 16192 10566 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 13035 16235 13093 16241
rect 13035 16232 13047 16235
rect 12584 16204 13047 16232
rect 12584 16192 12590 16204
rect 13035 16201 13047 16204
rect 13081 16201 13093 16235
rect 13035 16195 13093 16201
rect 13403 16235 13461 16241
rect 13403 16201 13415 16235
rect 13449 16232 13461 16235
rect 13538 16232 13544 16244
rect 13449 16204 13544 16232
rect 13449 16201 13461 16204
rect 13403 16195 13461 16201
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 15289 16235 15347 16241
rect 15289 16201 15301 16235
rect 15335 16232 15347 16235
rect 15378 16232 15384 16244
rect 15335 16204 15384 16232
rect 15335 16201 15347 16204
rect 15289 16195 15347 16201
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 16298 16192 16304 16244
rect 16356 16232 16362 16244
rect 17221 16235 17279 16241
rect 17221 16232 17233 16235
rect 16356 16204 17233 16232
rect 16356 16192 16362 16204
rect 17221 16201 17233 16204
rect 17267 16201 17279 16235
rect 17221 16195 17279 16201
rect 17681 16235 17739 16241
rect 17681 16201 17693 16235
rect 17727 16232 17739 16235
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 17727 16204 18061 16232
rect 17727 16201 17739 16204
rect 17681 16195 17739 16201
rect 18049 16201 18061 16204
rect 18095 16201 18107 16235
rect 18049 16195 18107 16201
rect 6270 16164 6276 16176
rect 3344 16136 6276 16164
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1688 15960 1716 16059
rect 2406 16056 2412 16108
rect 2464 16056 2470 16108
rect 2590 16056 2596 16108
rect 2648 16056 2654 16108
rect 3344 16105 3372 16136
rect 6270 16124 6276 16136
rect 6328 16124 6334 16176
rect 6730 16124 6736 16176
rect 6788 16124 6794 16176
rect 10965 16167 11023 16173
rect 10965 16133 10977 16167
rect 11011 16164 11023 16167
rect 13814 16164 13820 16176
rect 11011 16136 11744 16164
rect 11011 16133 11023 16136
rect 10965 16127 11023 16133
rect 11716 16108 11744 16136
rect 13372 16136 13820 16164
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16065 3387 16099
rect 3329 16059 3387 16065
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 3605 16099 3663 16105
rect 3605 16096 3617 16099
rect 3476 16068 3617 16096
rect 3476 16056 3482 16068
rect 3605 16065 3617 16068
rect 3651 16065 3663 16099
rect 3605 16059 3663 16065
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 4614 16096 4620 16108
rect 3835 16068 4620 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 5626 16056 5632 16108
rect 5684 16056 5690 16108
rect 7009 16099 7067 16105
rect 7009 16096 7021 16099
rect 6656 16068 7021 16096
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 2924 16000 3157 16028
rect 2924 15988 2930 16000
rect 3145 15997 3157 16000
rect 3191 16028 3203 16031
rect 3970 16028 3976 16040
rect 3191 16000 3976 16028
rect 3191 15997 3203 16000
rect 3145 15991 3203 15997
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 4154 15988 4160 16040
rect 4212 16028 4218 16040
rect 5350 16028 5356 16040
rect 4212 16000 5356 16028
rect 4212 15988 4218 16000
rect 5350 15988 5356 16000
rect 5408 16028 5414 16040
rect 5813 16031 5871 16037
rect 5813 16028 5825 16031
rect 5408 16000 5825 16028
rect 5408 15988 5414 16000
rect 5813 15997 5825 16000
rect 5859 15997 5871 16031
rect 5813 15991 5871 15997
rect 6365 16031 6423 16037
rect 6365 15997 6377 16031
rect 6411 16028 6423 16031
rect 6454 16028 6460 16040
rect 6411 16000 6460 16028
rect 6411 15997 6423 16000
rect 6365 15991 6423 15997
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 6086 15960 6092 15972
rect 1688 15932 6092 15960
rect 6086 15920 6092 15932
rect 6144 15920 6150 15972
rect 6178 15920 6184 15972
rect 6236 15960 6242 15972
rect 6549 15963 6607 15969
rect 6549 15960 6561 15963
rect 6236 15932 6561 15960
rect 6236 15920 6242 15932
rect 6549 15929 6561 15932
rect 6595 15929 6607 15963
rect 6549 15923 6607 15929
rect 842 15852 848 15904
rect 900 15892 906 15904
rect 1489 15895 1547 15901
rect 1489 15892 1501 15895
rect 900 15864 1501 15892
rect 900 15852 906 15864
rect 1489 15861 1501 15864
rect 1535 15861 1547 15895
rect 1489 15855 1547 15861
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15892 2835 15895
rect 4062 15892 4068 15904
rect 2823 15864 4068 15892
rect 2823 15861 2835 15864
rect 2777 15855 2835 15861
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 5261 15895 5319 15901
rect 5261 15861 5273 15895
rect 5307 15892 5319 15895
rect 5442 15892 5448 15904
rect 5307 15864 5448 15892
rect 5307 15861 5319 15864
rect 5261 15855 5319 15861
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 5902 15852 5908 15904
rect 5960 15892 5966 15904
rect 6457 15895 6515 15901
rect 6457 15892 6469 15895
rect 5960 15864 6469 15892
rect 5960 15852 5966 15864
rect 6457 15861 6469 15864
rect 6503 15892 6515 15895
rect 6656 15892 6684 16068
rect 7009 16065 7021 16068
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 8662 16056 8668 16108
rect 8720 16056 8726 16108
rect 10388 16099 10446 16105
rect 10388 16065 10400 16099
rect 10434 16096 10446 16099
rect 10870 16096 10876 16108
rect 10434 16068 10876 16096
rect 10434 16065 10446 16068
rect 10388 16059 10446 16065
rect 10870 16056 10876 16068
rect 10928 16056 10934 16108
rect 11698 16105 11704 16108
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16096 11115 16099
rect 11563 16099 11621 16105
rect 11563 16096 11575 16099
rect 11103 16068 11575 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 11563 16065 11575 16068
rect 11609 16065 11621 16099
rect 11563 16059 11621 16065
rect 11666 16099 11704 16105
rect 11666 16065 11678 16099
rect 11666 16059 11704 16065
rect 11698 16056 11704 16059
rect 11756 16056 11762 16108
rect 13138 16099 13196 16105
rect 13138 16065 13150 16099
rect 13184 16096 13196 16099
rect 13372 16096 13400 16136
rect 13814 16124 13820 16136
rect 13872 16164 13878 16176
rect 14550 16164 14556 16176
rect 13872 16136 14556 16164
rect 13872 16124 13878 16136
rect 14550 16124 14556 16136
rect 14608 16124 14614 16176
rect 13184 16068 13400 16096
rect 13184 16065 13196 16068
rect 13138 16059 13196 16065
rect 13446 16056 13452 16108
rect 13504 16105 13510 16108
rect 13504 16099 13532 16105
rect 13520 16065 13532 16099
rect 13504 16059 13532 16065
rect 13504 16056 13510 16059
rect 15654 16056 15660 16108
rect 15712 16056 15718 16108
rect 17589 16099 17647 16105
rect 17589 16065 17601 16099
rect 17635 16096 17647 16099
rect 18322 16096 18328 16108
rect 17635 16068 18328 16096
rect 17635 16065 17647 16068
rect 17589 16059 17647 16065
rect 18322 16056 18328 16068
rect 18380 16056 18386 16108
rect 18414 16056 18420 16108
rect 18472 16056 18478 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 18877 16099 18935 16105
rect 18877 16096 18889 16099
rect 18555 16068 18889 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 18877 16065 18889 16068
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 22002 16056 22008 16108
rect 22060 16056 22066 16108
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 11241 16031 11299 16037
rect 11241 16028 11253 16031
rect 10652 16000 11253 16028
rect 10652 15988 10658 16000
rect 11241 15997 11253 16000
rect 11287 16028 11299 16031
rect 12618 16028 12624 16040
rect 11287 16000 12624 16028
rect 11287 15997 11299 16000
rect 11241 15991 11299 15997
rect 12618 15988 12624 16000
rect 12676 15988 12682 16040
rect 15746 15988 15752 16040
rect 15804 15988 15810 16040
rect 15838 15988 15844 16040
rect 15896 16028 15902 16040
rect 17402 16028 17408 16040
rect 15896 16000 17408 16028
rect 15896 15988 15902 16000
rect 17402 15988 17408 16000
rect 17460 16028 17466 16040
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 17460 16000 17785 16028
rect 17460 15988 17466 16000
rect 17773 15997 17785 16000
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 18601 16031 18659 16037
rect 18601 15997 18613 16031
rect 18647 15997 18659 16031
rect 18601 15991 18659 15997
rect 8849 15963 8907 15969
rect 8849 15929 8861 15963
rect 8895 15960 8907 15963
rect 12158 15960 12164 15972
rect 8895 15932 12164 15960
rect 8895 15929 8907 15932
rect 8849 15923 8907 15929
rect 12158 15920 12164 15932
rect 12216 15920 12222 15972
rect 16298 15920 16304 15972
rect 16356 15960 16362 15972
rect 18616 15960 18644 15991
rect 18874 15960 18880 15972
rect 16356 15932 18880 15960
rect 16356 15920 16362 15932
rect 18874 15920 18880 15932
rect 18932 15920 18938 15972
rect 6503 15864 6684 15892
rect 6733 15895 6791 15901
rect 6503 15861 6515 15864
rect 6457 15855 6515 15861
rect 6733 15861 6745 15895
rect 6779 15892 6791 15895
rect 7466 15892 7472 15904
rect 6779 15864 7472 15892
rect 6779 15861 6791 15864
rect 6733 15855 6791 15861
rect 7466 15852 7472 15864
rect 7524 15852 7530 15904
rect 10502 15901 10508 15904
rect 10459 15895 10508 15901
rect 10459 15861 10471 15895
rect 10505 15861 10508 15895
rect 10459 15855 10508 15861
rect 10502 15852 10508 15855
rect 10560 15852 10566 15904
rect 16206 15852 16212 15904
rect 16264 15852 16270 15904
rect 21082 15852 21088 15904
rect 21140 15892 21146 15904
rect 21821 15895 21879 15901
rect 21821 15892 21833 15895
rect 21140 15864 21833 15892
rect 21140 15852 21146 15864
rect 21821 15861 21833 15864
rect 21867 15861 21879 15895
rect 21821 15855 21879 15861
rect 1104 15802 22356 15824
rect 1104 15750 3606 15802
rect 3658 15750 3670 15802
rect 3722 15750 3734 15802
rect 3786 15750 3798 15802
rect 3850 15750 3862 15802
rect 3914 15750 8919 15802
rect 8971 15750 8983 15802
rect 9035 15750 9047 15802
rect 9099 15750 9111 15802
rect 9163 15750 9175 15802
rect 9227 15750 14232 15802
rect 14284 15750 14296 15802
rect 14348 15750 14360 15802
rect 14412 15750 14424 15802
rect 14476 15750 14488 15802
rect 14540 15750 19545 15802
rect 19597 15750 19609 15802
rect 19661 15750 19673 15802
rect 19725 15750 19737 15802
rect 19789 15750 19801 15802
rect 19853 15750 22356 15802
rect 1104 15728 22356 15750
rect 2406 15648 2412 15700
rect 2464 15648 2470 15700
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 3237 15691 3295 15697
rect 3237 15688 3249 15691
rect 2648 15660 3249 15688
rect 2648 15648 2654 15660
rect 3237 15657 3249 15660
rect 3283 15657 3295 15691
rect 3237 15651 3295 15657
rect 5902 15648 5908 15700
rect 5960 15648 5966 15700
rect 6086 15648 6092 15700
rect 6144 15688 6150 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 6144 15660 6285 15688
rect 6144 15648 6150 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 6273 15651 6331 15657
rect 7742 15648 7748 15700
rect 7800 15648 7806 15700
rect 10505 15691 10563 15697
rect 10505 15657 10517 15691
rect 10551 15688 10563 15691
rect 10778 15688 10784 15700
rect 10551 15660 10784 15688
rect 10551 15657 10563 15660
rect 10505 15651 10563 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 12437 15691 12495 15697
rect 12437 15688 12449 15691
rect 11940 15660 12449 15688
rect 11940 15648 11946 15660
rect 12437 15657 12449 15660
rect 12483 15657 12495 15691
rect 12437 15651 12495 15657
rect 15746 15648 15752 15700
rect 15804 15648 15810 15700
rect 18414 15648 18420 15700
rect 18472 15648 18478 15700
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 19521 15691 19579 15697
rect 19521 15688 19533 15691
rect 19392 15660 19533 15688
rect 19392 15648 19398 15660
rect 19521 15657 19533 15660
rect 19567 15657 19579 15691
rect 19521 15651 19579 15657
rect 2866 15580 2872 15632
rect 2924 15580 2930 15632
rect 4154 15620 4160 15632
rect 3896 15592 4160 15620
rect 1762 15512 1768 15564
rect 1820 15552 1826 15564
rect 1857 15555 1915 15561
rect 1857 15552 1869 15555
rect 1820 15524 1869 15552
rect 1820 15512 1826 15524
rect 1857 15521 1869 15524
rect 1903 15552 1915 15555
rect 2130 15552 2136 15564
rect 1903 15524 2136 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 2130 15512 2136 15524
rect 2188 15512 2194 15564
rect 2685 15555 2743 15561
rect 2685 15521 2697 15555
rect 2731 15552 2743 15555
rect 2884 15552 2912 15580
rect 3896 15561 3924 15592
rect 4154 15580 4160 15592
rect 4212 15580 4218 15632
rect 5810 15620 5816 15632
rect 5368 15592 5816 15620
rect 2731 15524 2912 15552
rect 3881 15555 3939 15561
rect 2731 15521 2743 15524
rect 2685 15515 2743 15521
rect 3881 15521 3893 15555
rect 3927 15521 3939 15555
rect 3881 15515 3939 15521
rect 4062 15512 4068 15564
rect 4120 15512 4126 15564
rect 5368 15561 5396 15592
rect 5810 15580 5816 15592
rect 5868 15580 5874 15632
rect 8570 15620 8576 15632
rect 8404 15592 8576 15620
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15521 5411 15555
rect 5353 15515 5411 15521
rect 5442 15512 5448 15564
rect 5500 15512 5506 15564
rect 8404 15561 8432 15592
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 8389 15555 8447 15561
rect 5552 15524 8340 15552
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 2869 15487 2927 15493
rect 2869 15484 2881 15487
rect 1596 15456 2881 15484
rect 1596 15357 1624 15456
rect 2869 15453 2881 15456
rect 2915 15484 2927 15487
rect 3462 15487 3520 15493
rect 3462 15484 3474 15487
rect 2915 15456 3474 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 3462 15453 3474 15456
rect 3508 15453 3520 15487
rect 3462 15447 3520 15453
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 5552 15484 5580 15524
rect 4028 15456 5580 15484
rect 4028 15444 4034 15456
rect 6454 15444 6460 15496
rect 6512 15444 6518 15496
rect 2038 15376 2044 15428
rect 2096 15376 2102 15428
rect 2777 15419 2835 15425
rect 2777 15385 2789 15419
rect 2823 15416 2835 15419
rect 3375 15419 3433 15425
rect 3375 15416 3387 15419
rect 2823 15388 3387 15416
rect 2823 15385 2835 15388
rect 2777 15379 2835 15385
rect 3375 15385 3387 15388
rect 3421 15385 3433 15419
rect 5537 15419 5595 15425
rect 5537 15416 5549 15419
rect 3375 15379 3433 15385
rect 4540 15388 5549 15416
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 1946 15308 1952 15360
rect 2004 15308 2010 15360
rect 2130 15308 2136 15360
rect 2188 15348 2194 15360
rect 2866 15348 2872 15360
rect 2188 15320 2872 15348
rect 2188 15308 2194 15320
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 4154 15308 4160 15360
rect 4212 15308 4218 15360
rect 4540 15357 4568 15388
rect 5537 15385 5549 15388
rect 5583 15385 5595 15419
rect 5537 15379 5595 15385
rect 7742 15376 7748 15428
rect 7800 15416 7806 15428
rect 8205 15419 8263 15425
rect 8205 15416 8217 15419
rect 7800 15388 8217 15416
rect 7800 15376 7806 15388
rect 8205 15385 8217 15388
rect 8251 15385 8263 15419
rect 8312 15416 8340 15524
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 10502 15512 10508 15564
rect 10560 15552 10566 15564
rect 10965 15555 11023 15561
rect 10965 15552 10977 15555
rect 10560 15524 10977 15552
rect 10560 15512 10566 15524
rect 10965 15521 10977 15524
rect 11011 15521 11023 15555
rect 10965 15515 11023 15521
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15521 11115 15555
rect 11057 15515 11115 15521
rect 8570 15444 8576 15496
rect 8628 15444 8634 15496
rect 10870 15444 10876 15496
rect 10928 15444 10934 15496
rect 11072 15484 11100 15515
rect 16206 15512 16212 15564
rect 16264 15512 16270 15564
rect 16298 15512 16304 15564
rect 16356 15512 16362 15564
rect 18877 15555 18935 15561
rect 18877 15521 18889 15555
rect 18923 15552 18935 15555
rect 19150 15552 19156 15564
rect 18923 15524 19156 15552
rect 18923 15521 18935 15524
rect 18877 15515 18935 15521
rect 19150 15512 19156 15524
rect 19208 15552 19214 15564
rect 19208 15524 19380 15552
rect 19208 15512 19214 15524
rect 10980 15456 11100 15484
rect 12621 15487 12679 15493
rect 8312 15388 8616 15416
rect 8205 15379 8263 15385
rect 4525 15351 4583 15357
rect 4525 15317 4537 15351
rect 4571 15317 4583 15351
rect 4525 15311 4583 15317
rect 8113 15351 8171 15357
rect 8113 15317 8125 15351
rect 8159 15348 8171 15351
rect 8478 15348 8484 15360
rect 8159 15320 8484 15348
rect 8159 15317 8171 15320
rect 8113 15311 8171 15317
rect 8478 15308 8484 15320
rect 8536 15308 8542 15360
rect 8588 15348 8616 15388
rect 10502 15376 10508 15428
rect 10560 15416 10566 15428
rect 10686 15416 10692 15428
rect 10560 15388 10692 15416
rect 10560 15376 10566 15388
rect 10686 15376 10692 15388
rect 10744 15416 10750 15428
rect 10980 15416 11008 15456
rect 12621 15453 12633 15487
rect 12667 15484 12679 15487
rect 13630 15484 13636 15496
rect 12667 15456 13636 15484
rect 12667 15453 12679 15456
rect 12621 15447 12679 15453
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 18782 15444 18788 15496
rect 18840 15484 18846 15496
rect 19352 15493 19380 15524
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 18840 15456 19257 15484
rect 18840 15444 18846 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 19337 15487 19395 15493
rect 19337 15453 19349 15487
rect 19383 15453 19395 15487
rect 19337 15447 19395 15453
rect 20508 15487 20566 15493
rect 20508 15453 20520 15487
rect 20554 15484 20566 15487
rect 21082 15484 21088 15496
rect 20554 15456 21088 15484
rect 20554 15453 20566 15456
rect 20508 15447 20566 15453
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 10744 15388 11008 15416
rect 10744 15376 10750 15388
rect 10594 15348 10600 15360
rect 8588 15320 10600 15348
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 16114 15308 16120 15360
rect 16172 15308 16178 15360
rect 20579 15351 20637 15357
rect 20579 15317 20591 15351
rect 20625 15348 20637 15351
rect 21174 15348 21180 15360
rect 20625 15320 21180 15348
rect 20625 15317 20637 15320
rect 20579 15311 20637 15317
rect 21174 15308 21180 15320
rect 21232 15308 21238 15360
rect 21818 15308 21824 15360
rect 21876 15308 21882 15360
rect 1104 15258 22356 15280
rect 1104 15206 4266 15258
rect 4318 15206 4330 15258
rect 4382 15206 4394 15258
rect 4446 15206 4458 15258
rect 4510 15206 4522 15258
rect 4574 15206 9579 15258
rect 9631 15206 9643 15258
rect 9695 15206 9707 15258
rect 9759 15206 9771 15258
rect 9823 15206 9835 15258
rect 9887 15206 14892 15258
rect 14944 15206 14956 15258
rect 15008 15206 15020 15258
rect 15072 15206 15084 15258
rect 15136 15206 15148 15258
rect 15200 15206 20205 15258
rect 20257 15206 20269 15258
rect 20321 15206 20333 15258
rect 20385 15206 20397 15258
rect 20449 15206 20461 15258
rect 20513 15206 22356 15258
rect 1104 15184 22356 15206
rect 1946 15104 1952 15156
rect 2004 15144 2010 15156
rect 2087 15147 2145 15153
rect 2087 15144 2099 15147
rect 2004 15116 2099 15144
rect 2004 15104 2010 15116
rect 2087 15113 2099 15116
rect 2133 15113 2145 15147
rect 2087 15107 2145 15113
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 3418 15144 3424 15156
rect 2915 15116 3424 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 3973 15147 4031 15153
rect 3973 15113 3985 15147
rect 4019 15144 4031 15147
rect 4154 15144 4160 15156
rect 4019 15116 4160 15144
rect 4019 15113 4031 15116
rect 3973 15107 4031 15113
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 7742 15104 7748 15156
rect 7800 15104 7806 15156
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8570 15144 8576 15156
rect 8251 15116 8576 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 12989 15147 13047 15153
rect 12989 15113 13001 15147
rect 13035 15144 13047 15147
rect 13630 15144 13636 15156
rect 13035 15116 13636 15144
rect 13035 15113 13047 15116
rect 12989 15107 13047 15113
rect 13630 15104 13636 15116
rect 13688 15104 13694 15156
rect 18322 15104 18328 15156
rect 18380 15104 18386 15156
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15113 19947 15147
rect 19889 15107 19947 15113
rect 4433 15079 4491 15085
rect 2516 15048 3188 15076
rect 2038 15017 2044 15020
rect 2016 15011 2044 15017
rect 2016 14977 2028 15011
rect 2016 14971 2044 14977
rect 2038 14968 2044 14971
rect 2096 14968 2102 15020
rect 2406 14900 2412 14952
rect 2464 14940 2470 14952
rect 2516 14949 2544 15048
rect 2590 14968 2596 15020
rect 2648 15008 2654 15020
rect 3160 15017 3188 15048
rect 4433 15045 4445 15079
rect 4479 15076 4491 15079
rect 4614 15076 4620 15088
rect 4479 15048 4620 15076
rect 4479 15045 4491 15048
rect 4433 15039 4491 15045
rect 4614 15036 4620 15048
rect 4672 15036 4678 15088
rect 15838 15076 15844 15088
rect 12452 15048 15844 15076
rect 2685 15011 2743 15017
rect 2685 15008 2697 15011
rect 2648 14980 2697 15008
rect 2648 14968 2654 14980
rect 2685 14977 2697 14980
rect 2731 15008 2743 15011
rect 3145 15011 3203 15017
rect 2731 14980 3096 15008
rect 2731 14977 2743 14980
rect 2685 14971 2743 14977
rect 3068 14949 3096 14980
rect 3145 14977 3157 15011
rect 3191 14977 3203 15011
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 3145 14971 3203 14977
rect 3528 14980 4905 15008
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 2464 14912 2513 14940
rect 2464 14900 2470 14912
rect 2501 14909 2513 14912
rect 2547 14909 2559 14943
rect 2501 14903 2559 14909
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14909 3111 14943
rect 3053 14903 3111 14909
rect 3068 14804 3096 14903
rect 3160 14872 3188 14971
rect 3528 14949 3556 14980
rect 4893 14977 4905 14980
rect 4939 15008 4951 15011
rect 5261 15011 5319 15017
rect 4939 14980 5212 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14909 3571 14943
rect 3513 14903 3571 14909
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 3605 14875 3663 14881
rect 3605 14872 3617 14875
rect 3160 14844 3617 14872
rect 3605 14841 3617 14844
rect 3651 14841 3663 14875
rect 3605 14835 3663 14841
rect 3804 14804 3832 14903
rect 4706 14900 4712 14952
rect 4764 14940 4770 14952
rect 5184 14949 5212 14980
rect 5261 14977 5273 15011
rect 5307 14977 5319 15011
rect 5261 14971 5319 14977
rect 4985 14943 5043 14949
rect 4985 14940 4997 14943
rect 4764 14912 4997 14940
rect 4764 14900 4770 14912
rect 4985 14909 4997 14912
rect 5031 14909 5043 14943
rect 4985 14903 5043 14909
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 5000 14872 5028 14903
rect 5276 14872 5304 14971
rect 7466 14968 7472 15020
rect 7524 14968 7530 15020
rect 8110 14968 8116 15020
rect 8168 14968 8174 15020
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 15008 8999 15011
rect 9398 15008 9404 15020
rect 8987 14980 9404 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 9398 14968 9404 14980
rect 9456 14968 9462 15020
rect 5626 14900 5632 14952
rect 5684 14900 5690 14952
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 8352 14912 8708 14940
rect 8352 14900 8358 14912
rect 5000 14844 5304 14872
rect 8478 14832 8484 14884
rect 8536 14872 8542 14884
rect 8573 14875 8631 14881
rect 8573 14872 8585 14875
rect 8536 14844 8585 14872
rect 8536 14832 8542 14844
rect 8573 14841 8585 14844
rect 8619 14841 8631 14875
rect 8680 14872 8708 14912
rect 8754 14900 8760 14952
rect 8812 14940 8818 14952
rect 12452 14949 12480 15048
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 17865 15079 17923 15085
rect 17865 15045 17877 15079
rect 17911 15076 17923 15079
rect 18233 15079 18291 15085
rect 17911 15048 18184 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 15008 12679 15011
rect 12986 15008 12992 15020
rect 12667 14980 12992 15008
rect 12667 14977 12679 14980
rect 12621 14971 12679 14977
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 15008 15991 15011
rect 16482 15008 16488 15020
rect 15979 14980 16488 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16482 14968 16488 14980
rect 16540 14968 16546 15020
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 9033 14943 9091 14949
rect 9033 14940 9045 14943
rect 8812 14912 9045 14940
rect 8812 14900 8818 14912
rect 9033 14909 9045 14912
rect 9079 14909 9091 14943
rect 9033 14903 9091 14909
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14940 12587 14943
rect 13078 14940 13084 14952
rect 12575 14912 13084 14940
rect 12575 14909 12587 14912
rect 12529 14903 12587 14909
rect 9140 14872 9168 14903
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 15841 14943 15899 14949
rect 15841 14940 15853 14943
rect 15528 14912 15853 14940
rect 15528 14900 15534 14912
rect 15841 14909 15853 14912
rect 15887 14909 15899 14943
rect 15841 14903 15899 14909
rect 16114 14900 16120 14952
rect 16172 14940 16178 14952
rect 16301 14943 16359 14949
rect 16301 14940 16313 14943
rect 16172 14912 16313 14940
rect 16172 14900 16178 14912
rect 16301 14909 16313 14912
rect 16347 14909 16359 14943
rect 16301 14903 16359 14909
rect 8680 14844 9168 14872
rect 18064 14872 18092 14971
rect 18156 14940 18184 15048
rect 18233 15045 18245 15079
rect 18279 15076 18291 15079
rect 19426 15076 19432 15088
rect 18279 15048 19432 15076
rect 18279 15045 18291 15048
rect 18233 15039 18291 15045
rect 19426 15036 19432 15048
rect 19484 15076 19490 15088
rect 19904 15076 19932 15107
rect 21082 15104 21088 15156
rect 21140 15104 21146 15156
rect 21174 15104 21180 15156
rect 21232 15104 21238 15156
rect 19484 15048 19932 15076
rect 20257 15079 20315 15085
rect 19484 15036 19490 15048
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 15008 18751 15011
rect 19242 15008 19248 15020
rect 18739 14980 19248 15008
rect 18739 14977 18751 14980
rect 18693 14971 18751 14977
rect 19242 14968 19248 14980
rect 19300 14968 19306 15020
rect 19536 15017 19564 15048
rect 20257 15045 20269 15079
rect 20303 15076 20315 15079
rect 20714 15076 20720 15088
rect 20303 15048 20720 15076
rect 20303 15045 20315 15048
rect 20257 15039 20315 15045
rect 20714 15036 20720 15048
rect 20772 15076 20778 15088
rect 21818 15076 21824 15088
rect 20772 15048 21824 15076
rect 20772 15036 20778 15048
rect 21818 15036 21824 15048
rect 21876 15036 21882 15088
rect 19521 15011 19579 15017
rect 19521 14977 19533 15011
rect 19567 14977 19579 15011
rect 19521 14971 19579 14977
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 20530 15008 20536 15020
rect 20128 14980 20536 15008
rect 20128 14968 20134 14980
rect 18785 14943 18843 14949
rect 18785 14940 18797 14943
rect 18156 14912 18797 14940
rect 18785 14909 18797 14912
rect 18831 14909 18843 14943
rect 18785 14903 18843 14909
rect 18874 14900 18880 14952
rect 18932 14900 18938 14952
rect 19150 14900 19156 14952
rect 19208 14900 19214 14952
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 19628 14872 19656 14903
rect 20346 14900 20352 14952
rect 20404 14900 20410 14952
rect 20456 14949 20484 14980
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 20441 14943 20499 14949
rect 20441 14909 20453 14943
rect 20487 14909 20499 14943
rect 20441 14903 20499 14909
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 21269 14943 21327 14949
rect 21269 14940 21281 14943
rect 20680 14912 21281 14940
rect 20680 14900 20686 14912
rect 21269 14909 21281 14912
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 19886 14872 19892 14884
rect 18064 14844 19892 14872
rect 8573 14835 8631 14841
rect 19886 14832 19892 14844
rect 19944 14872 19950 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 19944 14844 20729 14872
rect 19944 14832 19950 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 20717 14835 20775 14841
rect 3068 14776 3832 14804
rect 7653 14807 7711 14813
rect 7653 14773 7665 14807
rect 7699 14804 7711 14807
rect 12894 14804 12900 14816
rect 7699 14776 12900 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 13449 14807 13507 14813
rect 13449 14773 13461 14807
rect 13495 14804 13507 14807
rect 13538 14804 13544 14816
rect 13495 14776 13544 14804
rect 13495 14773 13507 14776
rect 13449 14767 13507 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 1104 14714 22356 14736
rect 1104 14662 3606 14714
rect 3658 14662 3670 14714
rect 3722 14662 3734 14714
rect 3786 14662 3798 14714
rect 3850 14662 3862 14714
rect 3914 14662 8919 14714
rect 8971 14662 8983 14714
rect 9035 14662 9047 14714
rect 9099 14662 9111 14714
rect 9163 14662 9175 14714
rect 9227 14662 14232 14714
rect 14284 14662 14296 14714
rect 14348 14662 14360 14714
rect 14412 14662 14424 14714
rect 14476 14662 14488 14714
rect 14540 14662 19545 14714
rect 19597 14662 19609 14714
rect 19661 14662 19673 14714
rect 19725 14662 19737 14714
rect 19789 14662 19801 14714
rect 19853 14662 22356 14714
rect 1104 14640 22356 14662
rect 6089 14603 6147 14609
rect 6089 14569 6101 14603
rect 6135 14600 6147 14603
rect 6454 14600 6460 14612
rect 6135 14572 6460 14600
rect 6135 14569 6147 14572
rect 6089 14563 6147 14569
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8812 14572 8953 14600
rect 8812 14560 8818 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 9398 14560 9404 14612
rect 9456 14560 9462 14612
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 9548 14572 9812 14600
rect 9548 14560 9554 14572
rect 1670 14492 1676 14544
rect 1728 14532 1734 14544
rect 9674 14532 9680 14544
rect 1728 14504 9680 14532
rect 1728 14492 1734 14504
rect 9674 14492 9680 14504
rect 9732 14492 9738 14544
rect 9784 14541 9812 14572
rect 10134 14560 10140 14612
rect 10192 14560 10198 14612
rect 13078 14560 13084 14612
rect 13136 14560 13142 14612
rect 15378 14600 15384 14612
rect 13832 14572 15384 14600
rect 9769 14535 9827 14541
rect 9769 14501 9781 14535
rect 9815 14501 9827 14535
rect 9769 14495 9827 14501
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 10226 14532 10232 14544
rect 9916 14504 10232 14532
rect 9916 14492 9922 14504
rect 10226 14492 10232 14504
rect 10284 14492 10290 14544
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14464 5595 14467
rect 5810 14464 5816 14476
rect 5583 14436 5816 14464
rect 5583 14433 5595 14436
rect 5537 14427 5595 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 5920 14436 6745 14464
rect 842 14356 848 14408
rect 900 14396 906 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 900 14368 1409 14396
rect 900 14356 906 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 5920 14396 5948 14436
rect 6733 14433 6745 14436
rect 6779 14464 6791 14467
rect 8294 14464 8300 14476
rect 6779 14436 8300 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 9048 14436 10088 14464
rect 5408 14368 5948 14396
rect 5408 14356 5414 14368
rect 6086 14356 6092 14408
rect 6144 14396 6150 14408
rect 6144 14368 6316 14396
rect 6144 14356 6150 14368
rect 5629 14331 5687 14337
rect 5629 14297 5641 14331
rect 5675 14328 5687 14331
rect 6288 14328 6316 14368
rect 6546 14356 6552 14408
rect 6604 14356 6610 14408
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14396 6699 14399
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 6687 14368 7021 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 6564 14328 6592 14356
rect 9048 14328 9076 14436
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 9214 14396 9220 14408
rect 9171 14368 9220 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 9214 14356 9220 14368
rect 9272 14396 9278 14408
rect 9585 14399 9643 14405
rect 9585 14396 9597 14399
rect 9272 14368 9597 14396
rect 9272 14356 9278 14368
rect 9585 14365 9597 14368
rect 9631 14365 9643 14399
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 9585 14359 9643 14365
rect 9692 14368 9873 14396
rect 5675 14300 6224 14328
rect 6288 14300 9076 14328
rect 9309 14331 9367 14337
rect 5675 14297 5687 14300
rect 5629 14291 5687 14297
rect 1578 14220 1584 14272
rect 1636 14220 1642 14272
rect 5718 14220 5724 14272
rect 5776 14220 5782 14272
rect 6196 14269 6224 14300
rect 9309 14297 9321 14331
rect 9355 14328 9367 14331
rect 9490 14328 9496 14340
rect 9355 14300 9496 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 9490 14288 9496 14300
rect 9548 14288 9554 14340
rect 6181 14263 6239 14269
rect 6181 14229 6193 14263
rect 6227 14229 6239 14263
rect 6181 14223 6239 14229
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 6549 14263 6607 14269
rect 6549 14260 6561 14263
rect 6420 14232 6561 14260
rect 6420 14220 6426 14232
rect 6549 14229 6561 14232
rect 6595 14229 6607 14263
rect 6549 14223 6607 14229
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 9398 14260 9404 14272
rect 8720 14232 9404 14260
rect 8720 14220 8726 14232
rect 9398 14220 9404 14232
rect 9456 14260 9462 14272
rect 9692 14260 9720 14368
rect 9861 14365 9873 14368
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 10060 14328 10088 14436
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 13722 14424 13728 14476
rect 13780 14424 13786 14476
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 12492 14368 13001 14396
rect 12492 14356 12498 14368
rect 12989 14365 13001 14368
rect 13035 14396 13047 14399
rect 13740 14396 13768 14424
rect 13035 14368 13768 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 12621 14331 12679 14337
rect 12621 14328 12633 14331
rect 10060 14300 12633 14328
rect 12621 14297 12633 14300
rect 12667 14328 12679 14331
rect 13832 14328 13860 14572
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 15470 14560 15476 14612
rect 15528 14560 15534 14612
rect 15565 14603 15623 14609
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 15654 14600 15660 14612
rect 15611 14572 15660 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 16298 14600 16304 14612
rect 16132 14572 16304 14600
rect 15286 14532 15292 14544
rect 15120 14504 15292 14532
rect 14642 14356 14648 14408
rect 14700 14356 14706 14408
rect 15120 14405 15148 14504
rect 15286 14492 15292 14504
rect 15344 14532 15350 14544
rect 16022 14532 16028 14544
rect 15344 14504 16028 14532
rect 15344 14492 15350 14504
rect 16022 14492 16028 14504
rect 16080 14492 16086 14544
rect 16132 14473 16160 14572
rect 16298 14560 16304 14572
rect 16356 14560 16362 14612
rect 16482 14560 16488 14612
rect 16540 14560 16546 14612
rect 19242 14560 19248 14612
rect 19300 14560 19306 14612
rect 20346 14560 20352 14612
rect 20404 14609 20410 14612
rect 20404 14603 20453 14609
rect 20404 14569 20407 14603
rect 20441 14569 20453 14603
rect 20404 14563 20453 14569
rect 20404 14560 20410 14563
rect 17865 14535 17923 14541
rect 17865 14532 17877 14535
rect 16224 14504 17877 14532
rect 15197 14467 15255 14473
rect 15197 14433 15209 14467
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 12667 14300 13860 14328
rect 12667 14297 12679 14300
rect 12621 14291 12679 14297
rect 9456 14232 9720 14260
rect 9456 14220 9462 14232
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 13449 14263 13507 14269
rect 13449 14260 13461 14263
rect 13412 14232 13461 14260
rect 13412 14220 13418 14232
rect 13449 14229 13461 14232
rect 13495 14229 13507 14263
rect 13449 14223 13507 14229
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 14185 14263 14243 14269
rect 14185 14260 14197 14263
rect 13780 14232 14197 14260
rect 13780 14220 13786 14232
rect 14185 14229 14197 14232
rect 14231 14229 14243 14263
rect 15212 14260 15240 14427
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14396 15991 14399
rect 16224 14396 16252 14504
rect 17865 14501 17877 14504
rect 17911 14501 17923 14535
rect 17865 14495 17923 14501
rect 19426 14492 19432 14544
rect 19484 14532 19490 14544
rect 19613 14535 19671 14541
rect 19613 14532 19625 14535
rect 19484 14504 19625 14532
rect 19484 14492 19490 14504
rect 19613 14501 19625 14504
rect 19659 14501 19671 14535
rect 19613 14495 19671 14501
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 16356 14436 17509 14464
rect 16356 14424 16362 14436
rect 17497 14433 17509 14436
rect 17543 14433 17555 14467
rect 17497 14427 17555 14433
rect 15979 14368 16252 14396
rect 16945 14399 17003 14405
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16945 14365 16957 14399
rect 16991 14396 17003 14399
rect 17310 14396 17316 14408
rect 16991 14368 17316 14396
rect 16991 14365 17003 14368
rect 16945 14359 17003 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14392 17463 14399
rect 17512 14392 17540 14427
rect 17451 14365 17540 14392
rect 17405 14364 17540 14365
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14365 17739 14399
rect 17405 14359 17463 14364
rect 17681 14359 17739 14365
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 19334 14396 19340 14408
rect 18739 14368 19340 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 16025 14331 16083 14337
rect 16025 14297 16037 14331
rect 16071 14328 16083 14331
rect 17037 14331 17095 14337
rect 17037 14328 17049 14331
rect 16071 14300 17049 14328
rect 16071 14297 16083 14300
rect 16025 14291 16083 14297
rect 17037 14297 17049 14300
rect 17083 14297 17095 14331
rect 17037 14291 17095 14297
rect 17221 14331 17279 14337
rect 17221 14297 17233 14331
rect 17267 14328 17279 14331
rect 17696 14328 17724 14359
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 19886 14396 19892 14408
rect 19475 14368 19892 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 20498 14399 20556 14405
rect 20498 14365 20510 14399
rect 20544 14396 20556 14399
rect 20714 14396 20720 14408
rect 20544 14368 20720 14396
rect 20544 14365 20556 14368
rect 20498 14359 20556 14365
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 22002 14356 22008 14408
rect 22060 14356 22066 14408
rect 17267 14300 17724 14328
rect 17267 14297 17279 14300
rect 17221 14291 17279 14297
rect 15378 14260 15384 14272
rect 15212 14232 15384 14260
rect 14185 14223 14243 14229
rect 15378 14220 15384 14232
rect 15436 14260 15442 14272
rect 16666 14260 16672 14272
rect 15436 14232 16672 14260
rect 15436 14220 15442 14232
rect 16666 14220 16672 14232
rect 16724 14260 16730 14272
rect 17236 14260 17264 14291
rect 18874 14288 18880 14340
rect 18932 14288 18938 14340
rect 16724 14232 17264 14260
rect 16724 14220 16730 14232
rect 17310 14220 17316 14272
rect 17368 14260 17374 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 17368 14232 18521 14260
rect 17368 14220 17374 14232
rect 18509 14229 18521 14232
rect 18555 14229 18567 14263
rect 18509 14223 18567 14229
rect 20530 14220 20536 14272
rect 20588 14260 20594 14272
rect 21821 14263 21879 14269
rect 21821 14260 21833 14263
rect 20588 14232 21833 14260
rect 20588 14220 20594 14232
rect 21821 14229 21833 14232
rect 21867 14229 21879 14263
rect 21821 14223 21879 14229
rect 1104 14170 22356 14192
rect 1104 14118 4266 14170
rect 4318 14118 4330 14170
rect 4382 14118 4394 14170
rect 4446 14118 4458 14170
rect 4510 14118 4522 14170
rect 4574 14118 9579 14170
rect 9631 14118 9643 14170
rect 9695 14118 9707 14170
rect 9759 14118 9771 14170
rect 9823 14118 9835 14170
rect 9887 14118 14892 14170
rect 14944 14118 14956 14170
rect 15008 14118 15020 14170
rect 15072 14118 15084 14170
rect 15136 14118 15148 14170
rect 15200 14118 20205 14170
rect 20257 14118 20269 14170
rect 20321 14118 20333 14170
rect 20385 14118 20397 14170
rect 20449 14118 20461 14170
rect 20513 14118 22356 14170
rect 1104 14096 22356 14118
rect 1578 14016 1584 14068
rect 1636 14056 1642 14068
rect 1636 14028 6914 14056
rect 1636 14016 1642 14028
rect 4617 13991 4675 13997
rect 4617 13957 4629 13991
rect 4663 13988 4675 13991
rect 5445 13991 5503 13997
rect 5445 13988 5457 13991
rect 4663 13960 5457 13988
rect 4663 13957 4675 13960
rect 4617 13951 4675 13957
rect 5445 13957 5457 13960
rect 5491 13957 5503 13991
rect 6886 13988 6914 14028
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 9861 14059 9919 14065
rect 9861 14056 9873 14059
rect 9364 14028 9873 14056
rect 9364 14016 9370 14028
rect 9861 14025 9873 14028
rect 9907 14025 9919 14059
rect 9861 14019 9919 14025
rect 10226 14016 10232 14068
rect 10284 14016 10290 14068
rect 12986 14016 12992 14068
rect 13044 14016 13050 14068
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 16485 14059 16543 14065
rect 16485 14056 16497 14059
rect 14700 14028 16497 14056
rect 14700 14016 14706 14028
rect 16485 14025 16497 14028
rect 16531 14025 16543 14059
rect 16485 14019 16543 14025
rect 16666 14016 16672 14068
rect 16724 14016 16730 14068
rect 17310 14056 17316 14068
rect 16960 14028 17316 14056
rect 10042 13988 10048 14000
rect 6886 13960 10048 13988
rect 5445 13951 5503 13957
rect 10042 13948 10048 13960
rect 10100 13948 10106 14000
rect 10244 13988 10272 14016
rect 10244 13960 10916 13988
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 4706 13920 4712 13932
rect 4479 13892 4712 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 4801 13923 4859 13929
rect 4801 13889 4813 13923
rect 4847 13920 4859 13923
rect 4890 13920 4896 13932
rect 4847 13892 4896 13920
rect 4847 13889 4859 13892
rect 4801 13883 4859 13889
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13920 5043 13923
rect 5258 13920 5264 13932
rect 5031 13892 5264 13920
rect 5031 13889 5043 13892
rect 4985 13883 5043 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 5902 13880 5908 13932
rect 5960 13880 5966 13932
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6733 13923 6791 13929
rect 6733 13920 6745 13923
rect 6043 13892 6745 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6733 13889 6745 13892
rect 6779 13920 6791 13923
rect 8202 13920 8208 13932
rect 6779 13892 8208 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 8662 13880 8668 13932
rect 8720 13880 8726 13932
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13920 9183 13923
rect 9674 13920 9680 13932
rect 9171 13892 9680 13920
rect 9171 13889 9183 13892
rect 9125 13883 9183 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 10888 13929 10916 13960
rect 11514 13948 11520 14000
rect 11572 13988 11578 14000
rect 11977 13991 12035 13997
rect 11977 13988 11989 13991
rect 11572 13960 11989 13988
rect 11572 13948 11578 13960
rect 11977 13957 11989 13960
rect 12023 13988 12035 13991
rect 12342 13988 12348 14000
rect 12023 13960 12348 13988
rect 12023 13957 12035 13960
rect 11977 13951 12035 13957
rect 12342 13948 12348 13960
rect 12400 13948 12406 14000
rect 15657 13991 15715 13997
rect 15657 13957 15669 13991
rect 15703 13988 15715 13991
rect 16301 13991 16359 13997
rect 16301 13988 16313 13991
rect 15703 13960 16313 13988
rect 15703 13957 15715 13960
rect 15657 13951 15715 13957
rect 16301 13957 16313 13960
rect 16347 13957 16359 13991
rect 16301 13951 16359 13957
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 10735 13923 10793 13929
rect 10735 13920 10747 13923
rect 10367 13892 10747 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 10735 13889 10747 13892
rect 10781 13889 10793 13923
rect 10735 13883 10793 13889
rect 10838 13923 10916 13929
rect 10838 13889 10850 13923
rect 10884 13892 10916 13923
rect 11082 13923 11140 13929
rect 11082 13920 11094 13923
rect 10980 13892 11094 13920
rect 10884 13889 10896 13892
rect 10838 13883 10896 13889
rect 1670 13852 1676 13864
rect 1596 13824 1676 13852
rect 1596 13793 1624 13824
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 5276 13852 5304 13880
rect 6086 13852 6092 13864
rect 5276 13824 6092 13852
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 6362 13812 6368 13864
rect 6420 13812 6426 13864
rect 6641 13855 6699 13861
rect 6641 13821 6653 13855
rect 6687 13821 6699 13855
rect 6641 13815 6699 13821
rect 1581 13787 1639 13793
rect 1581 13753 1593 13787
rect 1627 13753 1639 13787
rect 1581 13747 1639 13753
rect 5902 13744 5908 13796
rect 5960 13784 5966 13796
rect 6656 13784 6684 13815
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 8168 13824 8309 13852
rect 8168 13812 8174 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13852 8815 13855
rect 9217 13855 9275 13861
rect 8803 13824 9168 13852
rect 8803 13821 8815 13824
rect 8757 13815 8815 13821
rect 5960 13756 6684 13784
rect 9140 13784 9168 13824
rect 9217 13821 9229 13855
rect 9263 13852 9275 13855
rect 9306 13852 9312 13864
rect 9263 13824 9312 13852
rect 9263 13821 9275 13824
rect 9217 13815 9275 13821
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 9416 13824 9505 13852
rect 9416 13784 9444 13824
rect 9493 13821 9505 13824
rect 9539 13852 9551 13855
rect 9950 13852 9956 13864
rect 9539 13824 9956 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10594 13852 10600 13864
rect 10551 13824 10600 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 9140 13756 9444 13784
rect 5960 13744 5966 13756
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10980 13784 11008 13892
rect 11082 13889 11094 13892
rect 11128 13889 11140 13923
rect 11082 13883 11140 13889
rect 11790 13880 11796 13932
rect 11848 13880 11854 13932
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 12529 13923 12587 13929
rect 12529 13920 12541 13923
rect 12207 13892 12541 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 12529 13889 12541 13892
rect 12575 13889 12587 13923
rect 12529 13883 12587 13889
rect 12618 13880 12624 13932
rect 12676 13880 12682 13932
rect 13722 13880 13728 13932
rect 13780 13880 13786 13932
rect 15378 13880 15384 13932
rect 15436 13880 15442 13932
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13920 15623 13923
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15611 13892 16129 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 12434 13812 12440 13864
rect 12492 13812 12498 13864
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13852 15255 13855
rect 15286 13852 15292 13864
rect 15243 13824 15292 13852
rect 15243 13821 15255 13824
rect 15197 13815 15255 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 15841 13855 15899 13861
rect 15841 13852 15853 13855
rect 15528 13824 15853 13852
rect 15528 13812 15534 13824
rect 15841 13821 15853 13824
rect 15887 13821 15899 13855
rect 15841 13815 15899 13821
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13852 16083 13855
rect 16960 13852 16988 14028
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18874 14056 18880 14068
rect 18647 14028 18880 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 21634 13988 21640 14000
rect 17083 13960 17724 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 17696 13929 17724 13960
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17543 13923 17601 13929
rect 17543 13920 17555 13923
rect 17175 13892 17555 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17543 13889 17555 13892
rect 17589 13889 17601 13923
rect 17543 13883 17601 13889
rect 17646 13923 17724 13929
rect 17646 13889 17658 13923
rect 17692 13920 17724 13923
rect 18708 13960 21640 13988
rect 18708 13920 18736 13960
rect 21634 13948 21640 13960
rect 21692 13948 21698 14000
rect 17692 13892 18736 13920
rect 18785 13923 18843 13929
rect 17692 13889 17704 13892
rect 17646 13883 17704 13889
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 19886 13920 19892 13932
rect 18831 13892 19892 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 19886 13880 19892 13892
rect 19944 13880 19950 13932
rect 22002 13880 22008 13932
rect 22060 13880 22066 13932
rect 16071 13824 16988 13852
rect 17221 13855 17279 13861
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 17221 13821 17233 13855
rect 17267 13821 17279 13855
rect 17221 13815 17279 13821
rect 18969 13855 19027 13861
rect 18969 13821 18981 13855
rect 19015 13852 19027 13855
rect 19426 13852 19432 13864
rect 19015 13824 19432 13852
rect 19015 13821 19027 13824
rect 18969 13815 19027 13821
rect 10100 13756 11008 13784
rect 10100 13744 10106 13756
rect 17126 13744 17132 13796
rect 17184 13784 17190 13796
rect 17236 13784 17264 13815
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20622 13784 20628 13796
rect 17184 13756 20628 13784
rect 17184 13744 17190 13756
rect 20622 13744 20628 13756
rect 20680 13744 20686 13796
rect 10318 13676 10324 13728
rect 10376 13716 10382 13728
rect 11011 13719 11069 13725
rect 11011 13716 11023 13719
rect 10376 13688 11023 13716
rect 10376 13676 10382 13688
rect 11011 13685 11023 13688
rect 11057 13685 11069 13719
rect 11011 13679 11069 13685
rect 21818 13676 21824 13728
rect 21876 13676 21882 13728
rect 1104 13626 22356 13648
rect 1104 13574 3606 13626
rect 3658 13574 3670 13626
rect 3722 13574 3734 13626
rect 3786 13574 3798 13626
rect 3850 13574 3862 13626
rect 3914 13574 8919 13626
rect 8971 13574 8983 13626
rect 9035 13574 9047 13626
rect 9099 13574 9111 13626
rect 9163 13574 9175 13626
rect 9227 13574 14232 13626
rect 14284 13574 14296 13626
rect 14348 13574 14360 13626
rect 14412 13574 14424 13626
rect 14476 13574 14488 13626
rect 14540 13574 19545 13626
rect 19597 13574 19609 13626
rect 19661 13574 19673 13626
rect 19725 13574 19737 13626
rect 19789 13574 19801 13626
rect 19853 13574 22356 13626
rect 1104 13552 22356 13574
rect 5350 13512 5356 13524
rect 4540 13484 5356 13512
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13345 4399 13379
rect 4540 13376 4568 13484
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 5445 13515 5503 13521
rect 5445 13481 5457 13515
rect 5491 13512 5503 13515
rect 5718 13512 5724 13524
rect 5491 13484 5724 13512
rect 5491 13481 5503 13484
rect 5445 13475 5503 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 9769 13515 9827 13521
rect 9769 13512 9781 13515
rect 8260 13484 9781 13512
rect 8260 13472 8266 13484
rect 9769 13481 9781 13484
rect 9815 13481 9827 13515
rect 9769 13475 9827 13481
rect 11333 13515 11391 13521
rect 11333 13481 11345 13515
rect 11379 13512 11391 13515
rect 12618 13512 12624 13524
rect 11379 13484 12624 13512
rect 11379 13481 11391 13484
rect 11333 13475 11391 13481
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 15286 13472 15292 13524
rect 15344 13472 15350 13524
rect 4617 13447 4675 13453
rect 4617 13413 4629 13447
rect 4663 13444 4675 13447
rect 5902 13444 5908 13456
rect 4663 13416 5908 13444
rect 4663 13413 4675 13416
rect 4617 13407 4675 13413
rect 5902 13404 5908 13416
rect 5960 13404 5966 13456
rect 8941 13447 8999 13453
rect 8941 13413 8953 13447
rect 8987 13444 8999 13447
rect 9674 13444 9680 13456
rect 8987 13416 9680 13444
rect 8987 13413 8999 13416
rect 8941 13407 8999 13413
rect 9674 13404 9680 13416
rect 9732 13444 9738 13456
rect 9861 13447 9919 13453
rect 9861 13444 9873 13447
rect 9732 13416 9873 13444
rect 9732 13404 9738 13416
rect 9861 13413 9873 13416
rect 9907 13413 9919 13447
rect 9861 13407 9919 13413
rect 11992 13416 15884 13444
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4540 13348 4813 13376
rect 4341 13339 4399 13345
rect 4801 13345 4813 13348
rect 4847 13345 4859 13379
rect 5074 13376 5080 13388
rect 4801 13339 4859 13345
rect 4908 13348 5080 13376
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 900 13280 1409 13308
rect 900 13268 906 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4356 13308 4384 13339
rect 4908 13308 4936 13348
rect 5074 13336 5080 13348
rect 5132 13376 5138 13388
rect 5132 13348 5764 13376
rect 5132 13336 5138 13348
rect 5736 13317 5764 13348
rect 5994 13336 6000 13388
rect 6052 13336 6058 13388
rect 9125 13379 9183 13385
rect 9125 13345 9137 13379
rect 9171 13376 9183 13379
rect 9306 13376 9312 13388
rect 9171 13348 9312 13376
rect 9171 13345 9183 13348
rect 9125 13339 9183 13345
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 10318 13336 10324 13388
rect 10376 13336 10382 13388
rect 10502 13336 10508 13388
rect 10560 13336 10566 13388
rect 11514 13336 11520 13388
rect 11572 13336 11578 13388
rect 11992 13385 12020 13416
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13345 12035 13379
rect 11977 13339 12035 13345
rect 4356 13280 4936 13308
rect 4985 13311 5043 13317
rect 4249 13271 4307 13277
rect 4985 13277 4997 13311
rect 5031 13308 5043 13311
rect 5537 13311 5595 13317
rect 5537 13308 5549 13311
rect 5031 13280 5549 13308
rect 5031 13277 5043 13280
rect 4985 13271 5043 13277
rect 5537 13277 5549 13280
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13308 5779 13311
rect 6181 13311 6239 13317
rect 6181 13308 6193 13311
rect 5767 13280 6193 13308
rect 5767 13277 5779 13280
rect 5721 13271 5779 13277
rect 6181 13277 6193 13280
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13308 9643 13311
rect 10134 13308 10140 13320
rect 9631 13280 10140 13308
rect 9631 13277 9643 13280
rect 9585 13271 9643 13277
rect 4264 13240 4292 13271
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 11716 13308 11744 13339
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12400 13348 12725 13376
rect 12400 13336 12406 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13345 13231 13379
rect 13173 13339 13231 13345
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13376 13967 13379
rect 14642 13376 14648 13388
rect 13955 13348 14648 13376
rect 13955 13345 13967 13348
rect 13909 13339 13967 13345
rect 11790 13308 11796 13320
rect 11716 13280 11796 13308
rect 11790 13268 11796 13280
rect 11848 13308 11854 13320
rect 12802 13308 12808 13320
rect 11848 13280 12808 13308
rect 11848 13268 11854 13280
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 13188 13308 13216 13339
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 15856 13385 15884 13416
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 20070 13376 20076 13388
rect 15887 13348 20076 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 20070 13336 20076 13348
rect 20128 13336 20134 13388
rect 13630 13308 13636 13320
rect 13188 13280 13636 13308
rect 13630 13268 13636 13280
rect 13688 13308 13694 13320
rect 13817 13311 13875 13317
rect 13817 13308 13829 13311
rect 13688 13280 13829 13308
rect 13688 13268 13694 13280
rect 13817 13277 13829 13280
rect 13863 13277 13875 13311
rect 13817 13271 13875 13277
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 16234 13311 16292 13317
rect 16234 13308 16246 13311
rect 15703 13280 16246 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 16234 13277 16246 13280
rect 16280 13308 16292 13311
rect 21726 13308 21732 13320
rect 16280 13280 21732 13308
rect 16280 13277 16292 13280
rect 16234 13271 16292 13277
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 22002 13268 22008 13320
rect 22060 13268 22066 13320
rect 4614 13240 4620 13252
rect 4264 13212 4620 13240
rect 4614 13200 4620 13212
rect 4672 13200 4678 13252
rect 5077 13243 5135 13249
rect 5077 13209 5089 13243
rect 5123 13240 5135 13243
rect 5123 13212 5672 13240
rect 5123 13209 5135 13212
rect 5077 13203 5135 13209
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 4154 13172 4160 13184
rect 1627 13144 4160 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 5644 13172 5672 13212
rect 5902 13200 5908 13252
rect 5960 13200 5966 13252
rect 9309 13243 9367 13249
rect 9309 13209 9321 13243
rect 9355 13240 9367 13243
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9355 13212 9413 13240
rect 9355 13209 9367 13212
rect 9309 13203 9367 13209
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9401 13203 9459 13209
rect 10042 13200 10048 13252
rect 10100 13240 10106 13252
rect 10229 13243 10287 13249
rect 10229 13240 10241 13243
rect 10100 13212 10241 13240
rect 10100 13200 10106 13212
rect 10229 13209 10241 13212
rect 10275 13209 10287 13243
rect 13078 13240 13084 13252
rect 10229 13203 10287 13209
rect 12176 13212 13084 13240
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 5644 13144 6377 13172
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 12066 13132 12072 13184
rect 12124 13132 12130 13184
rect 12176 13181 12204 13212
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 13354 13200 13360 13252
rect 13412 13200 13418 13252
rect 12161 13175 12219 13181
rect 12161 13141 12173 13175
rect 12207 13172 12219 13175
rect 12250 13172 12256 13184
rect 12207 13144 12256 13172
rect 12207 13141 12219 13144
rect 12161 13135 12219 13141
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12802 13172 12808 13184
rect 12575 13144 12808 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 15749 13175 15807 13181
rect 15749 13141 15761 13175
rect 15795 13172 15807 13175
rect 16163 13175 16221 13181
rect 16163 13172 16175 13175
rect 15795 13144 16175 13172
rect 15795 13141 15807 13144
rect 15749 13135 15807 13141
rect 16163 13141 16175 13144
rect 16209 13141 16221 13175
rect 16163 13135 16221 13141
rect 19610 13132 19616 13184
rect 19668 13172 19674 13184
rect 21821 13175 21879 13181
rect 21821 13172 21833 13175
rect 19668 13144 21833 13172
rect 19668 13132 19674 13144
rect 21821 13141 21833 13144
rect 21867 13141 21879 13175
rect 21821 13135 21879 13141
rect 1104 13082 22356 13104
rect 1104 13030 4266 13082
rect 4318 13030 4330 13082
rect 4382 13030 4394 13082
rect 4446 13030 4458 13082
rect 4510 13030 4522 13082
rect 4574 13030 9579 13082
rect 9631 13030 9643 13082
rect 9695 13030 9707 13082
rect 9759 13030 9771 13082
rect 9823 13030 9835 13082
rect 9887 13030 14892 13082
rect 14944 13030 14956 13082
rect 15008 13030 15020 13082
rect 15072 13030 15084 13082
rect 15136 13030 15148 13082
rect 15200 13030 20205 13082
rect 20257 13030 20269 13082
rect 20321 13030 20333 13082
rect 20385 13030 20397 13082
rect 20449 13030 20461 13082
rect 20513 13030 22356 13082
rect 1104 13008 22356 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 3881 12971 3939 12977
rect 1627 12940 2774 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 2746 12900 2774 12940
rect 3881 12937 3893 12971
rect 3927 12968 3939 12971
rect 4154 12968 4160 12980
rect 3927 12940 4160 12968
rect 3927 12937 3939 12940
rect 3881 12931 3939 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4249 12971 4307 12977
rect 4249 12937 4261 12971
rect 4295 12968 4307 12971
rect 4614 12968 4620 12980
rect 4295 12940 4620 12968
rect 4295 12937 4307 12940
rect 4249 12931 4307 12937
rect 4614 12928 4620 12940
rect 4672 12968 4678 12980
rect 4672 12940 4844 12968
rect 4672 12928 4678 12940
rect 4706 12900 4712 12912
rect 2746 12872 4712 12900
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 4816 12832 4844 12940
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 4948 12940 5181 12968
rect 4948 12928 4954 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 5169 12931 5227 12937
rect 12066 12928 12072 12980
rect 12124 12977 12130 12980
rect 12124 12971 12173 12977
rect 12124 12937 12127 12971
rect 12161 12937 12173 12971
rect 12124 12931 12173 12937
rect 12989 12971 13047 12977
rect 12989 12937 13001 12971
rect 13035 12937 13047 12971
rect 12989 12931 13047 12937
rect 12124 12928 12130 12931
rect 7300 12872 7972 12900
rect 5902 12832 5908 12844
rect 4816 12804 5908 12832
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 2924 12736 3617 12764
rect 2924 12724 2930 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12764 3847 12767
rect 4246 12764 4252 12776
rect 3835 12736 4252 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 4433 12767 4491 12773
rect 4433 12733 4445 12767
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 3142 12656 3148 12708
rect 3200 12696 3206 12708
rect 4448 12696 4476 12727
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 5552 12773 5580 12804
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7300 12841 7328 12872
rect 7944 12841 7972 12872
rect 12342 12860 12348 12912
rect 12400 12900 12406 12912
rect 13004 12900 13032 12931
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 21818 12968 21824 12980
rect 13136 12940 21824 12968
rect 13136 12928 13142 12940
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 12400 12872 13308 12900
rect 12400 12860 12406 12872
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 7248 12804 7297 12832
rect 7248 12792 7254 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12832 7435 12835
rect 7791 12835 7849 12841
rect 7791 12832 7803 12835
rect 7423 12804 7803 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7791 12801 7803 12804
rect 7837 12801 7849 12835
rect 7791 12795 7849 12801
rect 7894 12835 7972 12841
rect 7894 12801 7906 12835
rect 7940 12804 7972 12835
rect 12044 12835 12102 12841
rect 7940 12801 7952 12804
rect 7894 12795 7952 12801
rect 12044 12801 12056 12835
rect 12090 12832 12102 12835
rect 12250 12832 12256 12844
rect 12090 12804 12256 12832
rect 12090 12801 12102 12804
rect 12044 12795 12102 12801
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 12618 12792 12624 12844
rect 12676 12832 12682 12844
rect 13280 12841 13308 12872
rect 13354 12860 13360 12912
rect 13412 12900 13418 12912
rect 13817 12903 13875 12909
rect 13817 12900 13829 12903
rect 13412 12872 13829 12900
rect 13412 12860 13418 12872
rect 13817 12869 13829 12872
rect 13863 12869 13875 12903
rect 13817 12863 13875 12869
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 19610 12900 19616 12912
rect 19392 12872 19616 12900
rect 19392 12860 19398 12872
rect 19610 12860 19616 12872
rect 19668 12860 19674 12912
rect 20441 12903 20499 12909
rect 20441 12869 20453 12903
rect 20487 12900 20499 12903
rect 20530 12900 20536 12912
rect 20487 12872 20536 12900
rect 20487 12869 20499 12872
rect 20441 12863 20499 12869
rect 20530 12860 20536 12872
rect 20588 12860 20594 12912
rect 13265 12835 13323 12841
rect 12676 12804 13216 12832
rect 12676 12792 12682 12804
rect 5353 12767 5411 12773
rect 5353 12764 5365 12767
rect 5092 12736 5365 12764
rect 5092 12708 5120 12736
rect 5353 12733 5365 12736
rect 5399 12733 5411 12767
rect 5353 12727 5411 12733
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 7558 12724 7564 12776
rect 7616 12724 7622 12776
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 3200 12668 4476 12696
rect 3200 12656 3206 12668
rect 4448 12628 4476 12668
rect 5074 12656 5080 12708
rect 5132 12656 5138 12708
rect 7650 12696 7656 12708
rect 5184 12668 7656 12696
rect 5184 12628 5212 12668
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 12452 12696 12480 12727
rect 12526 12724 12532 12776
rect 12584 12724 12590 12776
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 12860 12736 13093 12764
rect 12860 12724 12866 12736
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13188 12764 13216 12804
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12832 13507 12835
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 13495 12804 13645 12832
rect 13495 12801 13507 12804
rect 13449 12795 13507 12801
rect 13633 12801 13645 12804
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 16546 12804 21864 12832
rect 16546 12764 16574 12804
rect 13188 12736 16574 12764
rect 13081 12727 13139 12733
rect 18230 12724 18236 12776
rect 18288 12764 18294 12776
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18288 12736 18705 12764
rect 18288 12724 18294 12736
rect 18693 12733 18705 12736
rect 18739 12764 18751 12767
rect 18739 12736 19380 12764
rect 18739 12733 18751 12736
rect 18693 12727 18751 12733
rect 15378 12696 15384 12708
rect 12452 12668 12940 12696
rect 4448 12600 5212 12628
rect 6914 12588 6920 12640
rect 6972 12588 6978 12640
rect 12912 12628 12940 12668
rect 13372 12668 15384 12696
rect 13372 12628 13400 12668
rect 15378 12656 15384 12668
rect 15436 12656 15442 12708
rect 18046 12656 18052 12708
rect 18104 12696 18110 12708
rect 18598 12696 18604 12708
rect 18104 12668 18604 12696
rect 18104 12656 18110 12668
rect 18598 12656 18604 12668
rect 18656 12696 18662 12708
rect 18877 12699 18935 12705
rect 18877 12696 18889 12699
rect 18656 12668 18889 12696
rect 18656 12656 18662 12668
rect 18877 12665 18889 12668
rect 18923 12696 18935 12699
rect 19245 12699 19303 12705
rect 19245 12696 19257 12699
rect 18923 12668 19257 12696
rect 18923 12665 18935 12668
rect 18877 12659 18935 12665
rect 19245 12665 19257 12668
rect 19291 12665 19303 12699
rect 19352 12696 19380 12736
rect 19426 12724 19432 12776
rect 19484 12764 19490 12776
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 19484 12736 19717 12764
rect 19484 12724 19490 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 19886 12724 19892 12776
rect 19944 12724 19950 12776
rect 20530 12724 20536 12776
rect 20588 12724 20594 12776
rect 20714 12724 20720 12776
rect 20772 12724 20778 12776
rect 21836 12705 21864 12804
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 20073 12699 20131 12705
rect 20073 12696 20085 12699
rect 19352 12668 20085 12696
rect 19245 12659 19303 12665
rect 20073 12665 20085 12668
rect 20119 12665 20131 12699
rect 20073 12659 20131 12665
rect 21821 12699 21879 12705
rect 21821 12665 21833 12699
rect 21867 12665 21879 12699
rect 21821 12659 21879 12665
rect 12912 12600 13400 12628
rect 14001 12631 14059 12637
rect 14001 12597 14013 12631
rect 14047 12628 14059 12631
rect 15286 12628 15292 12640
rect 14047 12600 15292 12628
rect 14047 12597 14059 12600
rect 14001 12591 14059 12597
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 18414 12588 18420 12640
rect 18472 12588 18478 12640
rect 18506 12588 18512 12640
rect 18564 12588 18570 12640
rect 1104 12538 22356 12560
rect 1104 12486 3606 12538
rect 3658 12486 3670 12538
rect 3722 12486 3734 12538
rect 3786 12486 3798 12538
rect 3850 12486 3862 12538
rect 3914 12486 8919 12538
rect 8971 12486 8983 12538
rect 9035 12486 9047 12538
rect 9099 12486 9111 12538
rect 9163 12486 9175 12538
rect 9227 12486 14232 12538
rect 14284 12486 14296 12538
rect 14348 12486 14360 12538
rect 14412 12486 14424 12538
rect 14476 12486 14488 12538
rect 14540 12486 19545 12538
rect 19597 12486 19609 12538
rect 19661 12486 19673 12538
rect 19725 12486 19737 12538
rect 19789 12486 19801 12538
rect 19853 12486 22356 12538
rect 1104 12464 22356 12486
rect 4246 12384 4252 12436
rect 4304 12433 4310 12436
rect 4304 12427 4353 12433
rect 4304 12393 4307 12427
rect 4341 12393 4353 12427
rect 4304 12387 4353 12393
rect 4304 12384 4310 12387
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 4755 12427 4813 12433
rect 4755 12424 4767 12427
rect 4672 12396 4767 12424
rect 4672 12384 4678 12396
rect 4755 12393 4767 12396
rect 4801 12393 4813 12427
rect 4755 12387 4813 12393
rect 9398 12384 9404 12436
rect 9456 12384 9462 12436
rect 12526 12384 12532 12436
rect 12584 12433 12590 12436
rect 12584 12427 12633 12433
rect 12584 12393 12587 12427
rect 12621 12393 12633 12427
rect 12584 12387 12633 12393
rect 12584 12384 12590 12387
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19567 12427 19625 12433
rect 19567 12424 19579 12427
rect 19484 12396 19579 12424
rect 19484 12384 19490 12396
rect 19567 12393 19579 12396
rect 19613 12393 19625 12427
rect 19567 12387 19625 12393
rect 19843 12427 19901 12433
rect 19843 12393 19855 12427
rect 19889 12424 19901 12427
rect 20530 12424 20536 12436
rect 19889 12396 20536 12424
rect 19889 12393 19901 12396
rect 19843 12387 19901 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 6549 12359 6607 12365
rect 6549 12325 6561 12359
rect 6595 12356 6607 12359
rect 6914 12356 6920 12368
rect 6595 12328 6920 12356
rect 6595 12325 6607 12328
rect 6549 12319 6607 12325
rect 6914 12316 6920 12328
rect 6972 12316 6978 12368
rect 14090 12316 14096 12368
rect 14148 12356 14154 12368
rect 14148 12328 19932 12356
rect 14148 12316 14154 12328
rect 19904 12300 19932 12328
rect 7650 12248 7656 12300
rect 7708 12288 7714 12300
rect 8110 12288 8116 12300
rect 7708 12260 8116 12288
rect 7708 12248 7714 12260
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10410 12288 10416 12300
rect 10367 12260 10416 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 17678 12288 17684 12300
rect 17451 12260 17684 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 17865 12291 17923 12297
rect 17865 12257 17877 12291
rect 17911 12288 17923 12291
rect 18230 12288 18236 12300
rect 17911 12260 18236 12288
rect 17911 12257 17923 12260
rect 17865 12251 17923 12257
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 18690 12248 18696 12300
rect 18748 12248 18754 12300
rect 19886 12248 19892 12300
rect 19944 12248 19950 12300
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4706 12229 4712 12232
rect 4366 12223 4424 12229
rect 4366 12220 4378 12223
rect 4212 12192 4378 12220
rect 4212 12180 4218 12192
rect 4366 12189 4378 12192
rect 4412 12189 4424 12223
rect 4366 12183 4424 12189
rect 4684 12223 4712 12229
rect 4684 12189 4696 12223
rect 4684 12183 4712 12189
rect 4706 12180 4712 12183
rect 4764 12180 4770 12232
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 7954 12223 8012 12229
rect 7954 12220 7966 12223
rect 6779 12192 7052 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 7024 12096 7052 12192
rect 7392 12192 7966 12220
rect 7392 12096 7420 12192
rect 7954 12189 7966 12192
rect 8000 12189 8012 12223
rect 7954 12183 8012 12189
rect 10134 12180 10140 12232
rect 10192 12180 10198 12232
rect 12618 12180 12624 12232
rect 12676 12229 12682 12232
rect 12676 12223 12704 12229
rect 12692 12189 12704 12223
rect 12676 12183 12704 12189
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 12676 12180 12682 12183
rect 8938 12112 8944 12164
rect 8996 12152 9002 12164
rect 9585 12155 9643 12161
rect 9585 12152 9597 12155
rect 8996 12124 9597 12152
rect 8996 12112 9002 12124
rect 9585 12121 9597 12124
rect 9631 12121 9643 12155
rect 9585 12115 9643 12121
rect 9769 12155 9827 12161
rect 9769 12121 9781 12155
rect 9815 12152 9827 12155
rect 9953 12155 10011 12161
rect 9953 12152 9965 12155
rect 9815 12124 9965 12152
rect 9815 12121 9827 12124
rect 9769 12115 9827 12121
rect 9953 12121 9965 12124
rect 9999 12121 10011 12155
rect 16868 12152 16896 12183
rect 17034 12180 17040 12232
rect 17092 12180 17098 12232
rect 17773 12223 17831 12229
rect 17773 12189 17785 12223
rect 17819 12220 17831 12223
rect 18046 12220 18052 12232
rect 17819 12192 18052 12220
rect 17819 12189 17831 12192
rect 17773 12183 17831 12189
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12220 18475 12223
rect 18506 12220 18512 12232
rect 18463 12192 18512 12220
rect 18463 12189 18475 12192
rect 18417 12183 18475 12189
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 19334 12180 19340 12232
rect 19392 12220 19398 12232
rect 19464 12223 19522 12229
rect 19464 12220 19476 12223
rect 19392 12192 19476 12220
rect 19392 12180 19398 12192
rect 19464 12189 19476 12192
rect 19510 12189 19522 12223
rect 19464 12183 19522 12189
rect 19772 12223 19830 12229
rect 19772 12189 19784 12223
rect 19818 12220 19830 12223
rect 20438 12220 20444 12232
rect 19818 12192 20444 12220
rect 19818 12189 19830 12192
rect 19772 12183 19830 12189
rect 20438 12180 20444 12192
rect 20496 12180 20502 12232
rect 17862 12152 17868 12164
rect 16868 12124 17868 12152
rect 9953 12115 10011 12121
rect 17862 12112 17868 12124
rect 17920 12112 17926 12164
rect 6914 12044 6920 12096
rect 6972 12044 6978 12096
rect 7006 12044 7012 12096
rect 7064 12044 7070 12096
rect 7374 12044 7380 12096
rect 7432 12044 7438 12096
rect 7469 12087 7527 12093
rect 7469 12053 7481 12087
rect 7515 12084 7527 12087
rect 7883 12087 7941 12093
rect 7883 12084 7895 12087
rect 7515 12056 7895 12084
rect 7515 12053 7527 12056
rect 7469 12047 7527 12053
rect 7883 12053 7895 12056
rect 7929 12053 7941 12087
rect 7883 12047 7941 12053
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17129 12087 17187 12093
rect 17129 12084 17141 12087
rect 17000 12056 17141 12084
rect 17000 12044 17006 12056
rect 17129 12053 17141 12056
rect 17175 12053 17187 12087
rect 17129 12047 17187 12053
rect 18046 12044 18052 12096
rect 18104 12044 18110 12096
rect 18322 12044 18328 12096
rect 18380 12084 18386 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 18380 12056 18521 12084
rect 18380 12044 18386 12056
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 18509 12047 18567 12053
rect 1104 11994 22356 12016
rect 1104 11942 4266 11994
rect 4318 11942 4330 11994
rect 4382 11942 4394 11994
rect 4446 11942 4458 11994
rect 4510 11942 4522 11994
rect 4574 11942 9579 11994
rect 9631 11942 9643 11994
rect 9695 11942 9707 11994
rect 9759 11942 9771 11994
rect 9823 11942 9835 11994
rect 9887 11942 14892 11994
rect 14944 11942 14956 11994
rect 15008 11942 15020 11994
rect 15072 11942 15084 11994
rect 15136 11942 15148 11994
rect 15200 11942 20205 11994
rect 20257 11942 20269 11994
rect 20321 11942 20333 11994
rect 20385 11942 20397 11994
rect 20449 11942 20461 11994
rect 20513 11942 22356 11994
rect 1104 11920 22356 11942
rect 6914 11840 6920 11892
rect 6972 11880 6978 11892
rect 7101 11883 7159 11889
rect 7101 11880 7113 11883
rect 6972 11852 7113 11880
rect 6972 11840 6978 11852
rect 7101 11849 7113 11852
rect 7147 11849 7159 11883
rect 7101 11843 7159 11849
rect 8938 11840 8944 11892
rect 8996 11840 9002 11892
rect 17129 11883 17187 11889
rect 17129 11849 17141 11883
rect 17175 11880 17187 11883
rect 17497 11883 17555 11889
rect 17497 11880 17509 11883
rect 17175 11852 17509 11880
rect 17175 11849 17187 11852
rect 17129 11843 17187 11849
rect 17497 11849 17509 11852
rect 17543 11849 17555 11883
rect 17497 11843 17555 11849
rect 17862 11840 17868 11892
rect 17920 11880 17926 11892
rect 17957 11883 18015 11889
rect 17957 11880 17969 11883
rect 17920 11852 17969 11880
rect 17920 11840 17926 11852
rect 17957 11849 17969 11852
rect 18003 11849 18015 11883
rect 17957 11843 18015 11849
rect 18322 11840 18328 11892
rect 18380 11840 18386 11892
rect 7193 11815 7251 11821
rect 7193 11781 7205 11815
rect 7239 11812 7251 11815
rect 8389 11815 8447 11821
rect 8389 11812 8401 11815
rect 7239 11784 8401 11812
rect 7239 11781 7251 11784
rect 7193 11775 7251 11781
rect 8389 11781 8401 11784
rect 8435 11781 8447 11815
rect 15749 11815 15807 11821
rect 8389 11775 8447 11781
rect 12544 11784 15700 11812
rect 842 11704 848 11756
rect 900 11744 906 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 900 11716 1409 11744
rect 900 11704 906 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1670 11704 1676 11756
rect 1728 11704 1734 11756
rect 1762 11704 1768 11756
rect 1820 11744 1826 11756
rect 2076 11747 2134 11753
rect 2076 11744 2088 11747
rect 1820 11716 2088 11744
rect 1820 11704 1826 11716
rect 2076 11713 2088 11716
rect 2122 11713 2134 11747
rect 2076 11707 2134 11713
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7745 11747 7803 11753
rect 7745 11744 7757 11747
rect 7064 11716 7757 11744
rect 7064 11704 7070 11716
rect 7745 11713 7757 11716
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 7190 11676 7196 11688
rect 1596 11648 7196 11676
rect 1596 11617 1624 11648
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7282 11636 7288 11688
rect 7340 11636 7346 11688
rect 7760 11676 7788 11707
rect 8018 11704 8024 11756
rect 8076 11704 8082 11756
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 8205 11707 8263 11713
rect 8588 11716 9229 11744
rect 8220 11676 8248 11707
rect 7760 11648 8248 11676
rect 8588 11620 8616 11716
rect 9217 11713 9229 11716
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11744 10287 11747
rect 10410 11744 10416 11756
rect 10275 11716 10416 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11388 11716 11529 11744
rect 11388 11704 11394 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 8803 11648 9137 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 9125 11645 9137 11648
rect 9171 11676 9183 11679
rect 9861 11679 9919 11685
rect 9861 11676 9873 11679
rect 9171 11648 9873 11676
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 9861 11645 9873 11648
rect 9907 11645 9919 11679
rect 9861 11639 9919 11645
rect 10134 11636 10140 11688
rect 10192 11676 10198 11688
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 10192 11648 10333 11676
rect 10192 11636 10198 11648
rect 10321 11645 10333 11648
rect 10367 11676 10379 11679
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10367 11648 10701 11676
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 10689 11645 10701 11648
rect 10735 11676 10747 11679
rect 10962 11676 10968 11688
rect 10735 11648 10968 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11577 1639 11611
rect 1581 11571 1639 11577
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 7374 11608 7380 11620
rect 1903 11580 7380 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 7929 11611 7987 11617
rect 7929 11608 7941 11611
rect 7484 11580 7941 11608
rect 2222 11549 2228 11552
rect 2179 11543 2228 11549
rect 2179 11509 2191 11543
rect 2225 11509 2228 11543
rect 2179 11503 2228 11509
rect 2222 11500 2228 11503
rect 2280 11500 2286 11552
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 6733 11543 6791 11549
rect 6733 11540 6745 11543
rect 6420 11512 6745 11540
rect 6420 11500 6426 11512
rect 6733 11509 6745 11512
rect 6779 11509 6791 11543
rect 6733 11503 6791 11509
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7484 11540 7512 11580
rect 7929 11577 7941 11580
rect 7975 11608 7987 11611
rect 8018 11608 8024 11620
rect 7975 11580 8024 11608
rect 7975 11577 7987 11580
rect 7929 11571 7987 11577
rect 8018 11568 8024 11580
rect 8076 11568 8082 11620
rect 8570 11568 8576 11620
rect 8628 11568 8634 11620
rect 10410 11568 10416 11620
rect 10468 11608 10474 11620
rect 10873 11611 10931 11617
rect 10873 11608 10885 11611
rect 10468 11580 10885 11608
rect 10468 11568 10474 11580
rect 10873 11577 10885 11580
rect 10919 11577 10931 11611
rect 10873 11571 10931 11577
rect 12544 11552 12572 11784
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 13872 11716 14289 11744
rect 13872 11704 13878 11716
rect 14277 11713 14289 11716
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15344 11716 15424 11744
rect 15344 11704 15350 11716
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 15396 11685 15424 11716
rect 14185 11679 14243 11685
rect 14185 11676 14197 11679
rect 14056 11648 14197 11676
rect 14056 11636 14062 11648
rect 14185 11645 14197 11648
rect 14231 11645 14243 11679
rect 14185 11639 14243 11645
rect 15381 11679 15439 11685
rect 15381 11645 15393 11679
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11645 15623 11679
rect 15672 11676 15700 11784
rect 15749 11781 15761 11815
rect 15795 11812 15807 11815
rect 16025 11815 16083 11821
rect 16025 11812 16037 11815
rect 15795 11784 16037 11812
rect 15795 11781 15807 11784
rect 15749 11775 15807 11781
rect 16025 11781 16037 11784
rect 16071 11781 16083 11815
rect 16025 11775 16083 11781
rect 17037 11815 17095 11821
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 18046 11812 18052 11824
rect 17083 11784 18052 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 18046 11772 18052 11784
rect 18104 11772 18110 11824
rect 18230 11772 18236 11824
rect 18288 11812 18294 11824
rect 18509 11815 18567 11821
rect 18509 11812 18521 11815
rect 18288 11784 18521 11812
rect 18288 11772 18294 11784
rect 18509 11781 18521 11784
rect 18555 11781 18567 11815
rect 18509 11775 18567 11781
rect 18598 11772 18604 11824
rect 18656 11812 18662 11824
rect 18693 11815 18751 11821
rect 18693 11812 18705 11815
rect 18656 11784 18705 11812
rect 18656 11772 18662 11784
rect 18693 11781 18705 11784
rect 18739 11781 18751 11815
rect 18693 11775 18751 11781
rect 15838 11704 15844 11756
rect 15896 11704 15902 11756
rect 15930 11704 15936 11756
rect 15988 11744 15994 11756
rect 17865 11747 17923 11753
rect 15988 11716 17356 11744
rect 15988 11704 15994 11716
rect 15672 11648 16896 11676
rect 15565 11639 15623 11645
rect 15580 11608 15608 11639
rect 14660 11580 15608 11608
rect 7156 11512 7512 11540
rect 7561 11543 7619 11549
rect 7156 11500 7162 11512
rect 7561 11509 7573 11543
rect 7607 11540 7619 11543
rect 7650 11540 7656 11552
rect 7607 11512 7656 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9456 11512 9597 11540
rect 9456 11500 9462 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 10594 11540 10600 11552
rect 10551 11512 10600 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 11701 11543 11759 11549
rect 11701 11509 11713 11543
rect 11747 11540 11759 11543
rect 12526 11540 12532 11552
rect 11747 11512 12532 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 14660 11549 14688 11580
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 14608 11512 14657 11540
rect 14608 11500 14614 11512
rect 14645 11509 14657 11512
rect 14691 11509 14703 11543
rect 14645 11503 14703 11509
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 14829 11543 14887 11549
rect 14829 11540 14841 11543
rect 14792 11512 14841 11540
rect 14792 11500 14798 11512
rect 14829 11509 14841 11512
rect 14875 11509 14887 11543
rect 14829 11503 14887 11509
rect 16206 11500 16212 11552
rect 16264 11500 16270 11552
rect 16666 11500 16672 11552
rect 16724 11500 16730 11552
rect 16868 11540 16896 11648
rect 16942 11636 16948 11688
rect 17000 11676 17006 11688
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 17000 11648 17233 11676
rect 17000 11636 17006 11648
rect 17221 11645 17233 11648
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 17328 11608 17356 11716
rect 17865 11713 17877 11747
rect 17911 11744 17923 11747
rect 18138 11744 18144 11756
rect 17911 11716 18144 11744
rect 17911 11713 17923 11716
rect 17865 11707 17923 11713
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 22002 11704 22008 11756
rect 22060 11704 22066 11756
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11676 18107 11679
rect 18690 11676 18696 11688
rect 18095 11648 18696 11676
rect 18095 11645 18107 11648
rect 18049 11639 18107 11645
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 21821 11611 21879 11617
rect 21821 11608 21833 11611
rect 17328 11580 21833 11608
rect 21821 11577 21833 11580
rect 21867 11577 21879 11611
rect 21821 11571 21879 11577
rect 20622 11540 20628 11552
rect 16868 11512 20628 11540
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 1104 11450 22356 11472
rect 1104 11398 3606 11450
rect 3658 11398 3670 11450
rect 3722 11398 3734 11450
rect 3786 11398 3798 11450
rect 3850 11398 3862 11450
rect 3914 11398 8919 11450
rect 8971 11398 8983 11450
rect 9035 11398 9047 11450
rect 9099 11398 9111 11450
rect 9163 11398 9175 11450
rect 9227 11398 14232 11450
rect 14284 11398 14296 11450
rect 14348 11398 14360 11450
rect 14412 11398 14424 11450
rect 14476 11398 14488 11450
rect 14540 11398 19545 11450
rect 19597 11398 19609 11450
rect 19661 11398 19673 11450
rect 19725 11398 19737 11450
rect 19789 11398 19801 11450
rect 19853 11398 22356 11450
rect 1104 11376 22356 11398
rect 8021 11339 8079 11345
rect 8021 11305 8033 11339
rect 8067 11336 8079 11339
rect 8570 11336 8576 11348
rect 8067 11308 8576 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 10468 11308 11989 11336
rect 10468 11296 10474 11308
rect 11977 11305 11989 11308
rect 12023 11305 12035 11339
rect 11977 11299 12035 11305
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 15838 11336 15844 11348
rect 13955 11308 15844 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 16960 11308 17540 11336
rect 2682 11228 2688 11280
rect 2740 11268 2746 11280
rect 2740 11240 10916 11268
rect 2740 11228 2746 11240
rect 1486 11092 1492 11144
rect 1544 11092 1550 11144
rect 2700 11141 2728 11228
rect 5258 11200 5264 11212
rect 3528 11172 5264 11200
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 3326 11132 3332 11144
rect 2915 11104 3332 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3528 11141 3556 11172
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 7006 11200 7012 11212
rect 6963 11172 7012 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 7190 11160 7196 11212
rect 7248 11160 7254 11212
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 7340 11172 9689 11200
rect 7340 11160 7346 11172
rect 9677 11169 9689 11172
rect 9723 11200 9735 11203
rect 10781 11203 10839 11209
rect 10781 11200 10793 11203
rect 9723 11172 10793 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 10781 11169 10793 11172
rect 10827 11169 10839 11203
rect 10888 11200 10916 11240
rect 10962 11228 10968 11280
rect 11020 11268 11026 11280
rect 11149 11271 11207 11277
rect 11149 11268 11161 11271
rect 11020 11240 11161 11268
rect 11020 11228 11026 11240
rect 11149 11237 11161 11240
rect 11195 11237 11207 11271
rect 11149 11231 11207 11237
rect 13464 11240 14504 11268
rect 11330 11200 11336 11212
rect 10888 11172 11336 11200
rect 10781 11163 10839 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 11790 11160 11796 11212
rect 11848 11160 11854 11212
rect 12526 11160 12532 11212
rect 12584 11160 12590 11212
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11101 3571 11135
rect 3513 11095 3571 11101
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11132 6883 11135
rect 7098 11132 7104 11144
rect 6871 11104 7104 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 7650 11092 7656 11144
rect 7708 11092 7714 11144
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9861 11135 9919 11141
rect 9861 11132 9873 11135
rect 9539 11104 9873 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9861 11101 9873 11104
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 13316 11135 13374 11141
rect 13316 11101 13328 11135
rect 13362 11132 13374 11135
rect 13464 11132 13492 11240
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 13630 11200 13636 11212
rect 13587 11172 13636 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11200 13783 11203
rect 13998 11200 14004 11212
rect 13771 11172 14004 11200
rect 13771 11169 13783 11172
rect 13725 11163 13783 11169
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 14090 11160 14096 11212
rect 14148 11200 14154 11212
rect 14185 11203 14243 11209
rect 14185 11200 14197 11203
rect 14148 11172 14197 11200
rect 14148 11160 14154 11172
rect 14185 11169 14197 11172
rect 14231 11169 14243 11203
rect 14185 11163 14243 11169
rect 14476 11141 14504 11240
rect 15378 11228 15384 11280
rect 15436 11268 15442 11280
rect 16482 11268 16488 11280
rect 15436 11240 16488 11268
rect 15436 11228 15442 11240
rect 15580 11209 15608 11240
rect 16482 11228 16488 11240
rect 16540 11228 16546 11280
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 15764 11172 16068 11200
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 13362 11104 13492 11132
rect 13648 11104 14381 11132
rect 13362 11101 13374 11104
rect 13316 11095 13374 11101
rect 1946 11024 1952 11076
rect 2004 11024 2010 11076
rect 3050 11024 3056 11076
rect 3108 11024 3114 11076
rect 3160 11036 3464 11064
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 1762 10996 1768 11008
rect 1719 10968 1768 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 1762 10956 1768 10968
rect 1820 10956 1826 11008
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 3160 10996 3188 11036
rect 3016 10968 3188 10996
rect 3016 10956 3022 10968
rect 3234 10956 3240 11008
rect 3292 10956 3298 11008
rect 3436 11005 3464 11036
rect 3970 11024 3976 11076
rect 4028 11064 4034 11076
rect 4525 11067 4583 11073
rect 4525 11064 4537 11067
rect 4028 11036 4537 11064
rect 4028 11024 4034 11036
rect 4525 11033 4537 11036
rect 4571 11033 4583 11067
rect 4525 11027 4583 11033
rect 4706 11024 4712 11076
rect 4764 11024 4770 11076
rect 4893 11067 4951 11073
rect 4893 11033 4905 11067
rect 4939 11064 4951 11067
rect 6730 11064 6736 11076
rect 4939 11036 6736 11064
rect 4939 11033 4951 11036
rect 4893 11027 4951 11033
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 7834 11024 7840 11076
rect 7892 11024 7898 11076
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 11790 11064 11796 11076
rect 8168 11036 11796 11064
rect 8168 11024 8174 11036
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 12437 11067 12495 11073
rect 12437 11064 12449 11067
rect 12124 11036 12449 11064
rect 12124 11024 12130 11036
rect 12437 11033 12449 11036
rect 12483 11033 12495 11067
rect 12437 11027 12495 11033
rect 13403 11067 13461 11073
rect 13403 11033 13415 11067
rect 13449 11064 13461 11067
rect 13648 11064 13676 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 15764 11132 15792 11172
rect 15930 11141 15936 11144
rect 14507 11104 15792 11132
rect 15898 11135 15936 11141
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 15898 11101 15910 11135
rect 15898 11095 15936 11101
rect 15930 11092 15936 11095
rect 15988 11092 15994 11144
rect 16040 11132 16068 11172
rect 16206 11160 16212 11212
rect 16264 11200 16270 11212
rect 16960 11209 16988 11308
rect 17405 11271 17463 11277
rect 17405 11237 17417 11271
rect 17451 11237 17463 11271
rect 17512 11268 17540 11308
rect 18138 11296 18144 11348
rect 18196 11296 18202 11348
rect 18233 11271 18291 11277
rect 18233 11268 18245 11271
rect 17512 11240 18245 11268
rect 17405 11231 17463 11237
rect 18233 11237 18245 11240
rect 18279 11237 18291 11271
rect 18233 11231 18291 11237
rect 21821 11271 21879 11277
rect 21821 11237 21833 11271
rect 21867 11237 21879 11271
rect 21821 11231 21879 11237
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 16264 11172 16957 11200
rect 16264 11160 16270 11172
rect 16945 11169 16957 11172
rect 16991 11169 17003 11203
rect 16945 11163 17003 11169
rect 17420 11132 17448 11231
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 17736 11172 18429 11200
rect 17736 11160 17742 11172
rect 18417 11169 18429 11172
rect 18463 11169 18475 11203
rect 21836 11200 21864 11231
rect 18417 11163 18475 11169
rect 18524 11172 21864 11200
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 16040 11104 16574 11132
rect 17420 11104 17785 11132
rect 13449 11036 13676 11064
rect 15289 11067 15347 11073
rect 13449 11033 13461 11036
rect 13403 11027 13461 11033
rect 15289 11033 15301 11067
rect 15335 11033 15347 11067
rect 15289 11027 15347 11033
rect 15381 11067 15439 11073
rect 15381 11033 15393 11067
rect 15427 11064 15439 11067
rect 15795 11067 15853 11073
rect 15795 11064 15807 11067
rect 15427 11036 15807 11064
rect 15427 11033 15439 11036
rect 15381 11027 15439 11033
rect 15795 11033 15807 11036
rect 15841 11033 15853 11067
rect 15795 11027 15853 11033
rect 3421 10999 3479 11005
rect 3421 10965 3433 10999
rect 3467 10996 3479 10999
rect 4062 10996 4068 11008
rect 3467 10968 4068 10996
rect 3467 10965 3479 10968
rect 3421 10959 3479 10965
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 9030 10956 9036 11008
rect 9088 10956 9094 11008
rect 10226 10956 10232 11008
rect 10284 10956 10290 11008
rect 10686 10956 10692 11008
rect 10744 10956 10750 11008
rect 11514 10956 11520 11008
rect 11572 10956 11578 11008
rect 11606 10956 11612 11008
rect 11664 10956 11670 11008
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 12345 10999 12403 11005
rect 12345 10996 12357 10999
rect 11940 10968 12357 10996
rect 11940 10956 11946 10968
rect 12345 10965 12357 10968
rect 12391 10965 12403 10999
rect 12345 10959 12403 10965
rect 14458 10956 14464 11008
rect 14516 10996 14522 11008
rect 14829 10999 14887 11005
rect 14829 10996 14841 10999
rect 14516 10968 14841 10996
rect 14516 10956 14522 10968
rect 14829 10965 14841 10968
rect 14875 10965 14887 10999
rect 14829 10959 14887 10965
rect 14921 10999 14979 11005
rect 14921 10965 14933 10999
rect 14967 10996 14979 10999
rect 15194 10996 15200 11008
rect 14967 10968 15200 10996
rect 14967 10965 14979 10968
rect 14921 10959 14979 10965
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15304 10996 15332 11027
rect 15948 10996 15976 11092
rect 16546 11064 16574 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 18524 11132 18552 11172
rect 17773 11095 17831 11101
rect 17880 11104 18552 11132
rect 18601 11135 18659 11141
rect 17880 11064 17908 11104
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 18647 11104 18889 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 18877 11101 18889 11104
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 22002 11092 22008 11144
rect 22060 11092 22066 11144
rect 16546 11036 17908 11064
rect 18506 11024 18512 11076
rect 18564 11064 18570 11076
rect 18693 11067 18751 11073
rect 18693 11064 18705 11067
rect 18564 11036 18705 11064
rect 18564 11024 18570 11036
rect 18693 11033 18705 11036
rect 18739 11033 18751 11067
rect 18693 11027 18751 11033
rect 15304 10968 15976 10996
rect 19058 10956 19064 11008
rect 19116 10956 19122 11008
rect 1104 10906 22356 10928
rect 1104 10854 4266 10906
rect 4318 10854 4330 10906
rect 4382 10854 4394 10906
rect 4446 10854 4458 10906
rect 4510 10854 4522 10906
rect 4574 10854 9579 10906
rect 9631 10854 9643 10906
rect 9695 10854 9707 10906
rect 9759 10854 9771 10906
rect 9823 10854 9835 10906
rect 9887 10854 14892 10906
rect 14944 10854 14956 10906
rect 15008 10854 15020 10906
rect 15072 10854 15084 10906
rect 15136 10854 15148 10906
rect 15200 10854 20205 10906
rect 20257 10854 20269 10906
rect 20321 10854 20333 10906
rect 20385 10854 20397 10906
rect 20449 10854 20461 10906
rect 20513 10854 22356 10906
rect 1104 10832 22356 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 3145 10795 3203 10801
rect 1627 10764 2774 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 2406 10684 2412 10736
rect 2464 10684 2470 10736
rect 2746 10724 2774 10764
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 3234 10792 3240 10804
rect 3191 10764 3240 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 5132 10764 5181 10792
rect 5132 10752 5138 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 9030 10752 9036 10804
rect 9088 10792 9094 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 9088 10764 9229 10792
rect 9088 10752 9094 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 9217 10755 9275 10761
rect 11606 10752 11612 10804
rect 11664 10801 11670 10804
rect 12066 10801 12072 10804
rect 11664 10795 11713 10801
rect 11664 10761 11667 10795
rect 11701 10761 11713 10795
rect 11664 10755 11713 10761
rect 12023 10795 12072 10801
rect 12023 10761 12035 10795
rect 12069 10761 12072 10795
rect 12023 10755 12072 10761
rect 11664 10752 11670 10755
rect 12066 10752 12072 10755
rect 12124 10752 12130 10804
rect 16482 10752 16488 10804
rect 16540 10792 16546 10804
rect 20714 10792 20720 10804
rect 16540 10764 20720 10792
rect 16540 10752 16546 10764
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 2746 10696 3280 10724
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 3142 10656 3148 10668
rect 1811 10628 2176 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 1949 10523 2007 10529
rect 1949 10489 1961 10523
rect 1995 10489 2007 10523
rect 2148 10520 2176 10628
rect 2240 10628 3148 10656
rect 2240 10597 2268 10628
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3252 10665 3280 10696
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 5905 10727 5963 10733
rect 5905 10724 5917 10727
rect 5868 10696 5917 10724
rect 5868 10684 5874 10696
rect 5905 10693 5917 10696
rect 5951 10693 5963 10727
rect 7374 10724 7380 10736
rect 5905 10687 5963 10693
rect 6656 10696 7380 10724
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 3384 10628 3893 10656
rect 3384 10616 3390 10628
rect 3881 10625 3893 10628
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4580 10628 5089 10656
rect 4580 10616 4586 10628
rect 5077 10625 5089 10628
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 2314 10548 2320 10600
rect 2372 10548 2378 10600
rect 2958 10548 2964 10600
rect 3016 10548 3022 10600
rect 3418 10548 3424 10600
rect 3476 10588 3482 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3476 10560 3801 10588
rect 3476 10548 3482 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 5353 10591 5411 10597
rect 5353 10588 5365 10591
rect 4120 10560 5365 10588
rect 4120 10548 4126 10560
rect 5353 10557 5365 10560
rect 5399 10588 5411 10591
rect 6656 10588 6684 10696
rect 7374 10684 7380 10696
rect 7432 10684 7438 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 7929 10727 7987 10733
rect 7929 10724 7941 10727
rect 7892 10696 7941 10724
rect 7892 10684 7898 10696
rect 7929 10693 7941 10696
rect 7975 10693 7987 10727
rect 7929 10687 7987 10693
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 10226 10724 10232 10736
rect 9171 10696 10232 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 11330 10684 11336 10736
rect 11388 10684 11394 10736
rect 15105 10727 15163 10733
rect 15105 10724 15117 10727
rect 14384 10696 15117 10724
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6788 10628 6929 10656
rect 6788 10616 6794 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 7190 10656 7196 10668
rect 6917 10619 6975 10625
rect 7024 10628 7196 10656
rect 5399 10560 6684 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 2777 10523 2835 10529
rect 2777 10520 2789 10523
rect 2148 10492 2789 10520
rect 1949 10483 2007 10489
rect 2777 10489 2789 10492
rect 2823 10520 2835 10523
rect 3050 10520 3056 10532
rect 2823 10492 3056 10520
rect 2823 10489 2835 10492
rect 2777 10483 2835 10489
rect 1964 10452 1992 10483
rect 3050 10480 3056 10492
rect 3108 10520 3114 10532
rect 3436 10520 3464 10548
rect 3108 10492 3464 10520
rect 3605 10523 3663 10529
rect 3108 10480 3114 10492
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 4982 10520 4988 10532
rect 3651 10492 4988 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 4982 10480 4988 10492
rect 5040 10480 5046 10532
rect 6932 10520 6960 10619
rect 7024 10597 7052 10628
rect 7190 10616 7196 10628
rect 7248 10656 7254 10668
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 7248 10628 7481 10656
rect 7248 10616 7254 10628
rect 7469 10625 7481 10628
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11726 10659 11784 10665
rect 11726 10656 11738 10659
rect 11664 10628 11738 10656
rect 11664 10616 11670 10628
rect 11726 10625 11738 10628
rect 11772 10625 11784 10659
rect 11726 10619 11784 10625
rect 11882 10616 11888 10668
rect 11940 10665 11946 10668
rect 11940 10659 11978 10665
rect 11966 10625 11978 10659
rect 11940 10619 11978 10625
rect 11940 10616 11946 10619
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 7392 10520 7420 10551
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14384 10588 14412 10696
rect 15105 10693 15117 10696
rect 15151 10724 15163 10727
rect 15286 10724 15292 10736
rect 15151 10696 15292 10724
rect 15151 10693 15163 10696
rect 15105 10687 15163 10693
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10656 14519 10659
rect 14734 10656 14740 10668
rect 14507 10628 14740 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10625 19303 10659
rect 19245 10619 19303 10625
rect 14056 10560 14412 10588
rect 14056 10548 14062 10560
rect 14550 10548 14556 10600
rect 14608 10548 14614 10600
rect 14936 10588 14964 10619
rect 14660 10560 14964 10588
rect 19260 10588 19288 10619
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 19392 10628 19441 10656
rect 19392 10616 19398 10628
rect 19429 10625 19441 10628
rect 19475 10656 19487 10659
rect 19889 10659 19947 10665
rect 19889 10656 19901 10659
rect 19475 10628 19901 10656
rect 19475 10625 19487 10628
rect 19429 10619 19487 10625
rect 19889 10625 19901 10628
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 20438 10616 20444 10668
rect 20496 10665 20502 10668
rect 20496 10659 20556 10665
rect 20496 10625 20510 10659
rect 20544 10656 20556 10659
rect 20544 10628 21864 10656
rect 20544 10625 20556 10628
rect 20496 10619 20556 10625
rect 20496 10616 20502 10619
rect 19705 10591 19763 10597
rect 19705 10588 19717 10591
rect 19260 10560 19717 10588
rect 6932 10492 7420 10520
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 7616 10492 10088 10520
rect 7616 10480 7622 10492
rect 3326 10452 3332 10464
rect 1964 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 4212 10424 4261 10452
rect 4212 10412 4218 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4249 10415 4307 10421
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 4890 10452 4896 10464
rect 4755 10424 4896 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5810 10412 5816 10464
rect 5868 10412 5874 10464
rect 7282 10412 7288 10464
rect 7340 10412 7346 10464
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 10060 10461 10088 10492
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 14458 10520 14464 10532
rect 13872 10492 14464 10520
rect 13872 10480 13878 10492
rect 14458 10480 14464 10492
rect 14516 10520 14522 10532
rect 14660 10520 14688 10560
rect 19705 10557 19717 10560
rect 19751 10557 19763 10591
rect 19705 10551 19763 10557
rect 14516 10492 14688 10520
rect 14829 10523 14887 10529
rect 14516 10480 14522 10492
rect 14829 10489 14841 10523
rect 14875 10520 14887 10523
rect 15470 10520 15476 10532
rect 14875 10492 15476 10520
rect 14875 10489 14887 10492
rect 14829 10483 14887 10489
rect 15470 10480 15476 10492
rect 15528 10480 15534 10532
rect 19720 10520 19748 10551
rect 19978 10520 19984 10532
rect 19720 10492 19984 10520
rect 19978 10480 19984 10492
rect 20036 10480 20042 10532
rect 21836 10529 21864 10628
rect 22002 10616 22008 10668
rect 22060 10616 22066 10668
rect 21821 10523 21879 10529
rect 21821 10489 21833 10523
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 8757 10455 8815 10461
rect 8757 10452 8769 10455
rect 8260 10424 8769 10452
rect 8260 10412 8266 10424
rect 8757 10421 8769 10424
rect 8803 10421 8815 10455
rect 8757 10415 8815 10421
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 11974 10452 11980 10464
rect 10091 10424 11980 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 11974 10412 11980 10424
rect 12032 10452 12038 10464
rect 14090 10452 14096 10464
rect 12032 10424 14096 10452
rect 12032 10412 12038 10424
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 14642 10452 14648 10464
rect 14231 10424 14648 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 15286 10412 15292 10464
rect 15344 10412 15350 10464
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19484 10424 19625 10452
rect 19484 10412 19490 10424
rect 19613 10421 19625 10424
rect 19659 10421 19671 10455
rect 19613 10415 19671 10421
rect 20070 10412 20076 10464
rect 20128 10412 20134 10464
rect 20395 10455 20453 10461
rect 20395 10421 20407 10455
rect 20441 10452 20453 10455
rect 20530 10452 20536 10464
rect 20441 10424 20536 10452
rect 20441 10421 20453 10424
rect 20395 10415 20453 10421
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 1104 10362 22356 10384
rect 1104 10310 3606 10362
rect 3658 10310 3670 10362
rect 3722 10310 3734 10362
rect 3786 10310 3798 10362
rect 3850 10310 3862 10362
rect 3914 10310 8919 10362
rect 8971 10310 8983 10362
rect 9035 10310 9047 10362
rect 9099 10310 9111 10362
rect 9163 10310 9175 10362
rect 9227 10310 14232 10362
rect 14284 10310 14296 10362
rect 14348 10310 14360 10362
rect 14412 10310 14424 10362
rect 14476 10310 14488 10362
rect 14540 10310 19545 10362
rect 19597 10310 19609 10362
rect 19661 10310 19673 10362
rect 19725 10310 19737 10362
rect 19789 10310 19801 10362
rect 19853 10310 22356 10362
rect 1104 10288 22356 10310
rect 2314 10208 2320 10260
rect 2372 10248 2378 10260
rect 2823 10251 2881 10257
rect 2823 10248 2835 10251
rect 2372 10220 2835 10248
rect 2372 10208 2378 10220
rect 2823 10217 2835 10220
rect 2869 10217 2881 10251
rect 2823 10211 2881 10217
rect 3421 10251 3479 10257
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 3970 10248 3976 10260
rect 3467 10220 3976 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4522 10208 4528 10260
rect 4580 10208 4586 10260
rect 5810 10248 5816 10260
rect 4908 10220 5816 10248
rect 2685 10183 2743 10189
rect 2685 10149 2697 10183
rect 2731 10149 2743 10183
rect 2685 10143 2743 10149
rect 3053 10183 3111 10189
rect 3053 10149 3065 10183
rect 3099 10180 3111 10183
rect 3326 10180 3332 10192
rect 3099 10152 3332 10180
rect 3099 10149 3111 10152
rect 3053 10143 3111 10149
rect 2130 10072 2136 10124
rect 2188 10072 2194 10124
rect 2222 10072 2228 10124
rect 2280 10072 2286 10124
rect 2700 10112 2728 10143
rect 3068 10112 3096 10143
rect 3326 10140 3332 10152
rect 3384 10140 3390 10192
rect 4154 10140 4160 10192
rect 4212 10140 4218 10192
rect 4908 10180 4936 10220
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 8168 10220 8309 10248
rect 8168 10208 8174 10220
rect 8297 10217 8309 10220
rect 8343 10217 8355 10251
rect 8297 10211 8355 10217
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 10781 10251 10839 10257
rect 10781 10248 10793 10251
rect 10744 10220 10793 10248
rect 10744 10208 10750 10220
rect 10781 10217 10793 10220
rect 10827 10217 10839 10251
rect 10781 10211 10839 10217
rect 12253 10251 12311 10257
rect 12253 10217 12265 10251
rect 12299 10248 12311 10251
rect 13170 10248 13176 10260
rect 12299 10220 13176 10248
rect 12299 10217 12311 10220
rect 12253 10211 12311 10217
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 18690 10248 18696 10260
rect 15436 10220 18696 10248
rect 15436 10208 15442 10220
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 19978 10248 19984 10260
rect 19576 10220 19984 10248
rect 19576 10208 19582 10220
rect 19978 10208 19984 10220
rect 20036 10248 20042 10260
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 20036 10220 20085 10248
rect 20036 10208 20042 10220
rect 20073 10217 20085 10220
rect 20119 10217 20131 10251
rect 20073 10211 20131 10217
rect 4816 10152 4936 10180
rect 5353 10183 5411 10189
rect 2700 10084 3096 10112
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3418 10112 3424 10124
rect 3283 10084 3424 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4172 10112 4200 10140
rect 4816 10121 4844 10152
rect 5353 10149 5365 10183
rect 5399 10149 5411 10183
rect 5353 10143 5411 10149
rect 12437 10183 12495 10189
rect 12437 10149 12449 10183
rect 12483 10149 12495 10183
rect 15562 10180 15568 10192
rect 12437 10143 12495 10149
rect 12636 10152 15568 10180
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 4172 10084 4261 10112
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 4249 10075 4307 10081
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 4890 10072 4896 10124
rect 4948 10072 4954 10124
rect 5368 10112 5396 10143
rect 7190 10112 7196 10124
rect 5368 10084 7196 10112
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 1688 9976 1716 10007
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 1820 10016 2329 10044
rect 1820 10004 1826 10016
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 2406 10004 2412 10056
rect 2464 10044 2470 10056
rect 2894 10047 2952 10053
rect 2894 10044 2906 10047
rect 2464 10016 2906 10044
rect 2464 10004 2470 10016
rect 2894 10013 2906 10016
rect 2940 10013 2952 10047
rect 2894 10007 2952 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4614 10044 4620 10056
rect 4203 10016 4620 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 4982 10004 4988 10056
rect 5040 10004 5046 10056
rect 5644 10053 5672 10084
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 12452 10112 12480 10143
rect 12084 10084 12480 10112
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 6730 10044 6736 10056
rect 6687 10016 6736 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10597 10047 10655 10053
rect 10597 10013 10609 10047
rect 10643 10044 10655 10047
rect 10962 10044 10968 10056
rect 10643 10016 10968 10044
rect 10643 10013 10655 10016
rect 10597 10007 10655 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 12084 10053 12112 10084
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 1688 9948 5488 9976
rect 1486 9868 1492 9920
rect 1544 9868 1550 9920
rect 5460 9917 5488 9948
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 7009 9979 7067 9985
rect 7009 9976 7021 9979
rect 6328 9948 7021 9976
rect 6328 9936 6334 9948
rect 7009 9945 7021 9948
rect 7055 9945 7067 9979
rect 12268 9976 12296 10007
rect 12342 10004 12348 10056
rect 12400 10004 12406 10056
rect 12548 10047 12606 10053
rect 12548 10013 12560 10047
rect 12594 10044 12606 10047
rect 12636 10044 12664 10152
rect 15562 10140 15568 10152
rect 15620 10140 15626 10192
rect 16669 10183 16727 10189
rect 16669 10149 16681 10183
rect 16715 10180 16727 10183
rect 21174 10180 21180 10192
rect 16715 10152 21180 10180
rect 16715 10149 16727 10152
rect 16669 10143 16727 10149
rect 21174 10140 21180 10152
rect 21232 10140 21238 10192
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10081 14519 10115
rect 14461 10075 14519 10081
rect 14553 10115 14611 10121
rect 14553 10081 14565 10115
rect 14599 10112 14611 10115
rect 15286 10112 15292 10124
rect 14599 10084 15292 10112
rect 14599 10081 14611 10084
rect 14553 10075 14611 10081
rect 12594 10016 12664 10044
rect 12594 10013 12606 10016
rect 12548 10007 12606 10013
rect 12710 10004 12716 10056
rect 12768 10004 12774 10056
rect 12802 10004 12808 10056
rect 12860 10004 12866 10056
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12952 10016 13185 10044
rect 12952 10004 12958 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 13081 9979 13139 9985
rect 12268 9948 12848 9976
rect 7009 9939 7067 9945
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9877 5503 9911
rect 5445 9871 5503 9877
rect 6454 9868 6460 9920
rect 6512 9868 6518 9920
rect 12434 9868 12440 9920
rect 12492 9868 12498 9920
rect 12820 9917 12848 9948
rect 13081 9945 13093 9979
rect 13127 9976 13139 9979
rect 13262 9976 13268 9988
rect 13127 9948 13268 9976
rect 13127 9945 13139 9948
rect 13081 9939 13139 9945
rect 13262 9936 13268 9948
rect 13320 9936 13326 9988
rect 14476 9976 14504 10075
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 16942 10072 16948 10124
rect 17000 10112 17006 10124
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 17000 10084 17417 10112
rect 17000 10072 17006 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10081 18383 10115
rect 18325 10075 18383 10081
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10044 16543 10047
rect 16666 10044 16672 10056
rect 16531 10016 16672 10044
rect 16531 10013 16543 10016
rect 16485 10007 16543 10013
rect 16666 10004 16672 10016
rect 16724 10044 16730 10056
rect 17862 10044 17868 10056
rect 16724 10016 17868 10044
rect 16724 10004 16730 10016
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 18340 10044 18368 10075
rect 18414 10072 18420 10124
rect 18472 10112 18478 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18472 10084 18521 10112
rect 18472 10072 18478 10084
rect 18509 10081 18521 10084
rect 18555 10112 18567 10115
rect 19058 10112 19064 10124
rect 18555 10084 19064 10112
rect 18555 10081 18567 10084
rect 18509 10075 18567 10081
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19484 10084 19717 10112
rect 19484 10072 19490 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 18690 10044 18696 10056
rect 18340 10016 18696 10044
rect 18690 10004 18696 10016
rect 18748 10044 18754 10056
rect 19812 10044 19840 10075
rect 20530 10072 20536 10124
rect 20588 10072 20594 10124
rect 20622 10072 20628 10124
rect 20680 10072 20686 10124
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 21453 10115 21511 10121
rect 21453 10112 21465 10115
rect 20772 10084 21465 10112
rect 20772 10072 20778 10084
rect 21453 10081 21465 10084
rect 21499 10081 21511 10115
rect 21453 10075 21511 10081
rect 18748 10016 19840 10044
rect 18748 10004 18754 10016
rect 20438 10004 20444 10056
rect 20496 10004 20502 10056
rect 21726 10004 21732 10056
rect 21784 10004 21790 10056
rect 15378 9976 15384 9988
rect 14476 9948 15384 9976
rect 15378 9936 15384 9948
rect 15436 9936 15442 9988
rect 17221 9979 17279 9985
rect 17221 9945 17233 9979
rect 17267 9976 17279 9979
rect 17267 9948 19288 9976
rect 17267 9945 17279 9948
rect 17221 9939 17279 9945
rect 12805 9911 12863 9917
rect 12805 9877 12817 9911
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 12989 9911 13047 9917
rect 12989 9877 13001 9911
rect 13035 9908 13047 9911
rect 14550 9908 14556 9920
rect 13035 9880 14556 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 14642 9868 14648 9920
rect 14700 9908 14706 9920
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14700 9880 15025 9908
rect 14700 9868 14706 9880
rect 15013 9877 15025 9880
rect 15059 9877 15071 9911
rect 15013 9871 15071 9877
rect 16850 9868 16856 9920
rect 16908 9868 16914 9920
rect 17313 9911 17371 9917
rect 17313 9877 17325 9911
rect 17359 9908 17371 9911
rect 17681 9911 17739 9917
rect 17681 9908 17693 9911
rect 17359 9880 17693 9908
rect 17359 9877 17371 9880
rect 17313 9871 17371 9877
rect 17681 9877 17693 9880
rect 17727 9877 17739 9911
rect 17681 9871 17739 9877
rect 18046 9868 18052 9920
rect 18104 9868 18110 9920
rect 18138 9868 18144 9920
rect 18196 9868 18202 9920
rect 18874 9868 18880 9920
rect 18932 9908 18938 9920
rect 19260 9917 19288 9948
rect 18969 9911 19027 9917
rect 18969 9908 18981 9911
rect 18932 9880 18981 9908
rect 18932 9868 18938 9880
rect 18969 9877 18981 9880
rect 19015 9877 19027 9911
rect 18969 9871 19027 9877
rect 19245 9911 19303 9917
rect 19245 9877 19257 9911
rect 19291 9877 19303 9911
rect 19245 9871 19303 9877
rect 19610 9868 19616 9920
rect 19668 9868 19674 9920
rect 20622 9868 20628 9920
rect 20680 9908 20686 9920
rect 20901 9911 20959 9917
rect 20901 9908 20913 9911
rect 20680 9880 20913 9908
rect 20680 9868 20686 9880
rect 20901 9877 20913 9880
rect 20947 9877 20959 9911
rect 20901 9871 20959 9877
rect 21266 9868 21272 9920
rect 21324 9868 21330 9920
rect 21358 9868 21364 9920
rect 21416 9868 21422 9920
rect 21910 9868 21916 9920
rect 21968 9868 21974 9920
rect 1104 9818 22356 9840
rect 1104 9766 4266 9818
rect 4318 9766 4330 9818
rect 4382 9766 4394 9818
rect 4446 9766 4458 9818
rect 4510 9766 4522 9818
rect 4574 9766 9579 9818
rect 9631 9766 9643 9818
rect 9695 9766 9707 9818
rect 9759 9766 9771 9818
rect 9823 9766 9835 9818
rect 9887 9766 14892 9818
rect 14944 9766 14956 9818
rect 15008 9766 15020 9818
rect 15072 9766 15084 9818
rect 15136 9766 15148 9818
rect 15200 9766 20205 9818
rect 20257 9766 20269 9818
rect 20321 9766 20333 9818
rect 20385 9766 20397 9818
rect 20449 9766 20461 9818
rect 20513 9766 22356 9818
rect 1104 9744 22356 9766
rect 2130 9664 2136 9716
rect 2188 9704 2194 9716
rect 7558 9704 7564 9716
rect 2188 9676 7564 9704
rect 2188 9664 2194 9676
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 16761 9707 16819 9713
rect 16761 9704 16773 9707
rect 12768 9676 16773 9704
rect 12768 9664 12774 9676
rect 16761 9673 16773 9676
rect 16807 9673 16819 9707
rect 16761 9667 16819 9673
rect 19610 9664 19616 9716
rect 19668 9704 19674 9716
rect 20625 9707 20683 9713
rect 20625 9704 20637 9707
rect 19668 9676 20637 9704
rect 19668 9664 19674 9676
rect 20625 9673 20637 9676
rect 20671 9673 20683 9707
rect 20625 9667 20683 9673
rect 20855 9707 20913 9713
rect 20855 9673 20867 9707
rect 20901 9704 20913 9707
rect 21358 9704 21364 9716
rect 20901 9676 21364 9704
rect 20901 9673 20913 9676
rect 20855 9667 20913 9673
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 4706 9596 4712 9648
rect 4764 9636 4770 9648
rect 4801 9639 4859 9645
rect 4801 9636 4813 9639
rect 4764 9608 4813 9636
rect 4764 9596 4770 9608
rect 4801 9605 4813 9608
rect 4847 9605 4859 9639
rect 4801 9599 4859 9605
rect 7837 9639 7895 9645
rect 7837 9605 7849 9639
rect 7883 9636 7895 9639
rect 12802 9636 12808 9648
rect 7883 9608 12808 9636
rect 7883 9605 7895 9608
rect 7837 9599 7895 9605
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 15197 9639 15255 9645
rect 15197 9605 15209 9639
rect 15243 9636 15255 9639
rect 15378 9636 15384 9648
rect 15243 9608 15384 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 16850 9636 16856 9648
rect 16316 9608 16856 9636
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4341 9571 4399 9577
rect 4341 9568 4353 9571
rect 4212 9540 4353 9568
rect 4212 9528 4218 9540
rect 4341 9537 4353 9540
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6730 9568 6736 9580
rect 6687 9540 6736 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 14734 9528 14740 9580
rect 14792 9568 14798 9580
rect 16316 9577 16344 9608
rect 16850 9596 16856 9608
rect 16908 9636 16914 9648
rect 16908 9608 17448 9636
rect 16908 9596 16914 9608
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14792 9540 15025 9568
rect 14792 9528 14798 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9537 16359 9571
rect 16301 9531 16359 9537
rect 16758 9528 16764 9580
rect 16816 9528 16822 9580
rect 17126 9528 17132 9580
rect 17184 9528 17190 9580
rect 17420 9577 17448 9608
rect 19260 9608 20116 9636
rect 17405 9571 17463 9577
rect 17405 9537 17417 9571
rect 17451 9537 17463 9571
rect 17405 9531 17463 9537
rect 17862 9528 17868 9580
rect 17920 9528 17926 9580
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 18196 9540 18245 9568
rect 18196 9528 18202 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 18874 9528 18880 9580
rect 18932 9528 18938 9580
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4172 9472 4261 9500
rect 4172 9444 4200 9472
rect 4249 9469 4261 9472
rect 4295 9500 4307 9503
rect 4614 9500 4620 9512
rect 4295 9472 4620 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 18104 9472 18521 9500
rect 18104 9460 18110 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 18782 9460 18788 9512
rect 18840 9500 18846 9512
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 18840 9472 19165 9500
rect 18840 9460 18846 9472
rect 19153 9469 19165 9472
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 4154 9392 4160 9444
rect 4212 9392 4218 9444
rect 16485 9435 16543 9441
rect 16485 9401 16497 9435
rect 16531 9432 16543 9435
rect 19260 9432 19288 9608
rect 19518 9528 19524 9580
rect 19576 9528 19582 9580
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 19981 9571 20039 9577
rect 19981 9568 19993 9571
rect 19944 9540 19993 9568
rect 19944 9528 19950 9540
rect 19981 9537 19993 9540
rect 20027 9537 20039 9571
rect 20088 9568 20116 9608
rect 20162 9596 20168 9648
rect 20220 9596 20226 9648
rect 21726 9636 21732 9648
rect 20272 9608 21732 9636
rect 20272 9568 20300 9608
rect 21726 9596 21732 9608
rect 21784 9596 21790 9648
rect 20088 9540 20300 9568
rect 20784 9571 20842 9577
rect 19981 9531 20039 9537
rect 20784 9537 20796 9571
rect 20830 9568 20842 9571
rect 21266 9568 21272 9580
rect 20830 9540 21272 9568
rect 20830 9537 20842 9540
rect 20784 9531 20842 9537
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 19392 9472 19441 9500
rect 19392 9460 19398 9472
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19536 9500 19564 9528
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 19536 9472 20269 9500
rect 19429 9463 19487 9469
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 20441 9503 20499 9509
rect 20441 9469 20453 9503
rect 20487 9500 20499 9503
rect 20622 9500 20628 9512
rect 20487 9472 20628 9500
rect 20487 9469 20499 9472
rect 20441 9463 20499 9469
rect 16531 9404 19288 9432
rect 19444 9432 19472 9463
rect 20456 9432 20484 9463
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 19444 9404 20484 9432
rect 16531 9401 16543 9404
rect 16485 9395 16543 9401
rect 15473 9367 15531 9373
rect 15473 9333 15485 9367
rect 15519 9364 15531 9367
rect 15562 9364 15568 9376
rect 15519 9336 15568 9364
rect 15519 9333 15531 9336
rect 15473 9327 15531 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 19797 9367 19855 9373
rect 19797 9333 19809 9367
rect 19843 9364 19855 9367
rect 19978 9364 19984 9376
rect 19843 9336 19984 9364
rect 19843 9333 19855 9336
rect 19797 9327 19855 9333
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 1104 9274 22356 9296
rect 1104 9222 3606 9274
rect 3658 9222 3670 9274
rect 3722 9222 3734 9274
rect 3786 9222 3798 9274
rect 3850 9222 3862 9274
rect 3914 9222 8919 9274
rect 8971 9222 8983 9274
rect 9035 9222 9047 9274
rect 9099 9222 9111 9274
rect 9163 9222 9175 9274
rect 9227 9222 14232 9274
rect 14284 9222 14296 9274
rect 14348 9222 14360 9274
rect 14412 9222 14424 9274
rect 14476 9222 14488 9274
rect 14540 9222 19545 9274
rect 19597 9222 19609 9274
rect 19661 9222 19673 9274
rect 19725 9222 19737 9274
rect 19789 9222 19801 9274
rect 19853 9222 22356 9274
rect 1104 9200 22356 9222
rect 6454 9160 6460 9172
rect 2746 9132 6460 9160
rect 842 9052 848 9104
rect 900 9092 906 9104
rect 1489 9095 1547 9101
rect 1489 9092 1501 9095
rect 900 9064 1501 9092
rect 900 9052 906 9064
rect 1489 9061 1501 9064
rect 1535 9061 1547 9095
rect 1489 9055 1547 9061
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 2746 8956 2774 9132
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 6730 9120 6736 9172
rect 6788 9120 6794 9172
rect 18785 9163 18843 9169
rect 18785 9129 18797 9163
rect 18831 9160 18843 9163
rect 19886 9160 19892 9172
rect 18831 9132 19892 9160
rect 18831 9129 18843 9132
rect 18785 9123 18843 9129
rect 19886 9120 19892 9132
rect 19944 9120 19950 9172
rect 7653 9095 7711 9101
rect 7653 9092 7665 9095
rect 1719 8928 2774 8956
rect 5184 9064 7665 9092
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 5184 8820 5212 9064
rect 7653 9061 7665 9064
rect 7699 9061 7711 9095
rect 7653 9055 7711 9061
rect 9398 9052 9404 9104
rect 9456 9092 9462 9104
rect 15013 9095 15071 9101
rect 9456 9064 12434 9092
rect 9456 9052 9462 9064
rect 5810 8984 5816 9036
rect 5868 9024 5874 9036
rect 6181 9027 6239 9033
rect 6181 9024 6193 9027
rect 5868 8996 6193 9024
rect 5868 8984 5874 8996
rect 6181 8993 6193 8996
rect 6227 9024 6239 9027
rect 6227 8996 7144 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 6273 8891 6331 8897
rect 6273 8857 6285 8891
rect 6319 8888 6331 8891
rect 7116 8888 7144 8996
rect 7374 8984 7380 9036
rect 7432 8984 7438 9036
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 7282 8956 7288 8968
rect 7239 8928 7288 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 9416 8965 9444 9052
rect 11514 9024 11520 9036
rect 9600 8996 11520 9024
rect 9600 8965 9628 8996
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 12406 9024 12434 9064
rect 15013 9061 15025 9095
rect 15059 9092 15071 9095
rect 15286 9092 15292 9104
rect 15059 9064 15292 9092
rect 15059 9061 15071 9064
rect 15013 9055 15071 9061
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 15436 9064 15700 9092
rect 15436 9052 15442 9064
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 12406 8996 14381 9024
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7800 8928 7849 8956
rect 7800 8916 7806 8928
rect 7837 8925 7849 8928
rect 7883 8956 7895 8959
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 7883 8928 8953 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 9416 8888 9444 8919
rect 6319 8860 6868 8888
rect 7116 8860 9444 8888
rect 6319 8857 6331 8860
rect 6273 8851 6331 8857
rect 6840 8829 6868 8860
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 9692 8888 9720 8919
rect 10318 8916 10324 8968
rect 10376 8965 10382 8968
rect 10376 8959 10414 8965
rect 10402 8925 10414 8959
rect 10376 8919 10414 8925
rect 10376 8916 10382 8919
rect 11054 8916 11060 8968
rect 11112 8916 11118 8968
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 9548 8860 9720 8888
rect 9548 8848 9554 8860
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 11256 8888 11284 8919
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 11834 8959 11892 8965
rect 11834 8956 11846 8959
rect 11388 8928 11846 8956
rect 11388 8916 11394 8928
rect 11834 8925 11846 8928
rect 11880 8925 11892 8959
rect 11834 8919 11892 8925
rect 12526 8916 12532 8968
rect 12584 8916 12590 8968
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8956 12679 8959
rect 12710 8956 12716 8968
rect 12667 8928 12716 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 12820 8965 12848 8996
rect 14369 8993 14381 8996
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 14476 8996 15332 9024
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 13354 8916 13360 8968
rect 13412 8916 13418 8968
rect 11747 8891 11805 8897
rect 11747 8888 11759 8891
rect 11256 8860 11759 8888
rect 11747 8857 11759 8860
rect 11793 8857 11805 8891
rect 11747 8851 11805 8857
rect 13265 8891 13323 8897
rect 13265 8857 13277 8891
rect 13311 8888 13323 8891
rect 14476 8888 14504 8996
rect 14642 8916 14648 8968
rect 14700 8916 14706 8968
rect 13311 8860 14504 8888
rect 14553 8891 14611 8897
rect 13311 8857 13323 8860
rect 13265 8851 13323 8857
rect 14553 8857 14565 8891
rect 14599 8888 14611 8891
rect 15304 8888 15332 8996
rect 15562 8984 15568 9036
rect 15620 8984 15626 9036
rect 15672 9033 15700 9064
rect 18414 9052 18420 9104
rect 18472 9052 18478 9104
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 8993 15715 9027
rect 16758 9024 16764 9036
rect 15657 8987 15715 8993
rect 15948 8996 16764 9024
rect 15470 8916 15476 8968
rect 15528 8916 15534 8968
rect 15948 8965 15976 8996
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 9024 18659 9027
rect 18782 9024 18788 9036
rect 18647 8996 18788 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8925 15991 8959
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 15933 8919 15991 8925
rect 16132 8928 21741 8956
rect 15948 8888 15976 8919
rect 14599 8860 15148 8888
rect 15304 8860 15976 8888
rect 14599 8857 14611 8860
rect 14553 8851 14611 8857
rect 1728 8792 5212 8820
rect 6825 8823 6883 8829
rect 1728 8780 1734 8792
rect 6825 8789 6837 8823
rect 6871 8789 6883 8823
rect 6825 8783 6883 8789
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 6972 8792 7297 8820
rect 6972 8780 6978 8792
rect 7285 8789 7297 8792
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 10410 8780 10416 8832
rect 10468 8829 10474 8832
rect 15120 8829 15148 8860
rect 16132 8829 16160 8928
rect 21729 8925 21741 8928
rect 21775 8925 21787 8959
rect 21729 8919 21787 8925
rect 10468 8823 10517 8829
rect 10468 8789 10471 8823
rect 10505 8789 10517 8823
rect 10468 8783 10517 8789
rect 15105 8823 15163 8829
rect 15105 8789 15117 8823
rect 15151 8789 15163 8823
rect 15105 8783 15163 8789
rect 16117 8823 16175 8829
rect 16117 8789 16129 8823
rect 16163 8789 16175 8823
rect 16117 8783 16175 8789
rect 10468 8780 10474 8783
rect 21910 8780 21916 8832
rect 21968 8780 21974 8832
rect 1104 8730 22356 8752
rect 1104 8678 4266 8730
rect 4318 8678 4330 8730
rect 4382 8678 4394 8730
rect 4446 8678 4458 8730
rect 4510 8678 4522 8730
rect 4574 8678 9579 8730
rect 9631 8678 9643 8730
rect 9695 8678 9707 8730
rect 9759 8678 9771 8730
rect 9823 8678 9835 8730
rect 9887 8678 14892 8730
rect 14944 8678 14956 8730
rect 15008 8678 15020 8730
rect 15072 8678 15084 8730
rect 15136 8678 15148 8730
rect 15200 8678 20205 8730
rect 20257 8678 20269 8730
rect 20321 8678 20333 8730
rect 20385 8678 20397 8730
rect 20449 8678 20461 8730
rect 20513 8678 22356 8730
rect 1104 8656 22356 8678
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4212 8588 4445 8616
rect 4212 8576 4218 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 8389 8619 8447 8625
rect 8389 8585 8401 8619
rect 8435 8616 8447 8619
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8435 8588 9229 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9217 8579 9275 8585
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9548 8588 9597 8616
rect 9548 8576 9554 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 3145 8551 3203 8557
rect 3145 8517 3157 8551
rect 3191 8548 3203 8551
rect 4338 8548 4344 8560
rect 3191 8520 4344 8548
rect 3191 8517 3203 8520
rect 3145 8511 3203 8517
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 10226 8548 10232 8560
rect 9048 8520 10232 8548
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3050 8480 3056 8492
rect 3007 8452 3056 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 2792 8412 2820 8443
rect 3050 8440 3056 8452
rect 3108 8480 3114 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3108 8452 3433 8480
rect 3108 8440 3114 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 4062 8440 4068 8492
rect 4120 8440 4126 8492
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 4212 8452 4261 8480
rect 4212 8440 4218 8452
rect 4249 8449 4261 8452
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 2792 8384 3280 8412
rect 3252 8356 3280 8384
rect 4706 8372 4712 8424
rect 4764 8372 4770 8424
rect 9048 8421 9076 8520
rect 10226 8508 10232 8520
rect 10284 8548 10290 8560
rect 10284 8520 10732 8548
rect 10284 8508 10290 8520
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9640 8452 9781 8480
rect 9640 8440 9646 8452
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 10594 8480 10600 8492
rect 10442 8466 10600 8480
rect 9769 8443 9827 8449
rect 10428 8452 10600 8466
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 9306 8412 9312 8424
rect 9171 8384 9312 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 3234 8304 3240 8356
rect 3292 8304 3298 8356
rect 3605 8347 3663 8353
rect 3605 8313 3617 8347
rect 3651 8344 3663 8347
rect 4246 8344 4252 8356
rect 3651 8316 4252 8344
rect 3651 8313 3663 8316
rect 3605 8307 3663 8313
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8344 5227 8347
rect 5534 8344 5540 8356
rect 5215 8316 5540 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 7098 8304 7104 8356
rect 7156 8344 7162 8356
rect 8021 8347 8079 8353
rect 8021 8344 8033 8347
rect 7156 8316 8033 8344
rect 7156 8304 7162 8316
rect 8021 8313 8033 8316
rect 8067 8313 8079 8347
rect 8021 8307 8079 8313
rect 5626 8236 5632 8288
rect 5684 8236 5690 8288
rect 8588 8276 8616 8375
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 10428 8412 10456 8452
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 10704 8480 10732 8520
rect 11514 8508 11520 8560
rect 11572 8508 11578 8560
rect 12710 8508 12716 8560
rect 12768 8508 12774 8560
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 10704 8452 11989 8480
rect 11977 8449 11989 8452
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8480 12219 8483
rect 12618 8480 12624 8492
rect 12207 8452 12624 8480
rect 12207 8449 12219 8452
rect 12161 8443 12219 8449
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13262 8480 13268 8492
rect 13219 8452 13268 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8480 14703 8483
rect 15286 8480 15292 8492
rect 14691 8452 15292 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8480 16727 8483
rect 17126 8480 17132 8492
rect 16715 8452 17132 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 19978 8480 19984 8492
rect 19352 8452 19984 8480
rect 9456 8384 10456 8412
rect 10781 8415 10839 8421
rect 9456 8372 9462 8384
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11238 8412 11244 8424
rect 10827 8384 11244 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 12250 8372 12256 8424
rect 12308 8372 12314 8424
rect 12636 8412 12664 8440
rect 13449 8415 13507 8421
rect 13449 8412 13461 8415
rect 12636 8384 13461 8412
rect 13449 8381 13461 8384
rect 13495 8381 13507 8415
rect 13449 8375 13507 8381
rect 19153 8415 19211 8421
rect 19153 8381 19165 8415
rect 19199 8412 19211 8415
rect 19242 8412 19248 8424
rect 19199 8384 19248 8412
rect 19199 8381 19211 8384
rect 19153 8375 19211 8381
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 19352 8421 19380 8452
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 19337 8415 19395 8421
rect 19337 8381 19349 8415
rect 19383 8381 19395 8415
rect 19337 8375 19395 8381
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8344 8815 8347
rect 9582 8344 9588 8356
rect 8803 8316 9588 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8344 14887 8347
rect 16206 8344 16212 8356
rect 14875 8316 16212 8344
rect 14875 8313 14887 8316
rect 14829 8307 14887 8313
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8344 16911 8347
rect 21376 8344 21404 8443
rect 16899 8316 21404 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 21542 8304 21548 8356
rect 21600 8304 21606 8356
rect 9398 8276 9404 8288
rect 8588 8248 9404 8276
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 17586 8236 17592 8288
rect 17644 8236 17650 8288
rect 18966 8236 18972 8288
rect 19024 8236 19030 8288
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 19521 8279 19579 8285
rect 19521 8276 19533 8279
rect 19484 8248 19533 8276
rect 19484 8236 19490 8248
rect 19521 8245 19533 8248
rect 19567 8245 19579 8279
rect 19521 8239 19579 8245
rect 1104 8186 22356 8208
rect 1104 8134 3606 8186
rect 3658 8134 3670 8186
rect 3722 8134 3734 8186
rect 3786 8134 3798 8186
rect 3850 8134 3862 8186
rect 3914 8134 8919 8186
rect 8971 8134 8983 8186
rect 9035 8134 9047 8186
rect 9099 8134 9111 8186
rect 9163 8134 9175 8186
rect 9227 8134 14232 8186
rect 14284 8134 14296 8186
rect 14348 8134 14360 8186
rect 14412 8134 14424 8186
rect 14476 8134 14488 8186
rect 14540 8134 19545 8186
rect 19597 8134 19609 8186
rect 19661 8134 19673 8186
rect 19725 8134 19737 8186
rect 19789 8134 19801 8186
rect 19853 8134 22356 8186
rect 1104 8112 22356 8134
rect 3050 8032 3056 8084
rect 3108 8032 3114 8084
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 4062 8072 4068 8084
rect 3559 8044 4068 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 9306 8072 9312 8084
rect 9171 8044 9312 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 11701 8075 11759 8081
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 12250 8072 12256 8084
rect 11747 8044 12256 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12584 8044 12633 8072
rect 12584 8032 12590 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 2225 8007 2283 8013
rect 2225 7973 2237 8007
rect 2271 8004 2283 8007
rect 3068 8004 3096 8032
rect 5442 8004 5448 8016
rect 2271 7976 3004 8004
rect 3068 7976 3372 8004
rect 2271 7973 2283 7976
rect 2225 7967 2283 7973
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 1946 7936 1952 7948
rect 1719 7908 1952 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 2976 7936 3004 7976
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 2547 7908 2774 7936
rect 2976 7908 3157 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 2746 7800 2774 7908
rect 3145 7905 3157 7908
rect 3191 7936 3203 7939
rect 3234 7936 3240 7948
rect 3191 7908 3240 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 3344 7945 3372 7976
rect 3988 7976 5448 8004
rect 3988 7945 4016 7976
rect 5442 7964 5448 7976
rect 5500 8004 5506 8016
rect 8205 8007 8263 8013
rect 5500 7976 5764 8004
rect 5500 7964 5506 7976
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7905 3387 7939
rect 3329 7899 3387 7905
rect 3973 7939 4031 7945
rect 3973 7905 3985 7939
rect 4019 7905 4031 7939
rect 3973 7899 4031 7905
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4338 7936 4344 7948
rect 4111 7908 4344 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 5626 7896 5632 7948
rect 5684 7896 5690 7948
rect 5736 7945 5764 7976
rect 8205 7973 8217 8007
rect 8251 8004 8263 8007
rect 12434 8004 12440 8016
rect 8251 7976 12440 8004
rect 8251 7973 8263 7976
rect 8205 7967 8263 7973
rect 12434 7964 12440 7976
rect 12492 7964 12498 8016
rect 15841 8007 15899 8013
rect 15841 7973 15853 8007
rect 15887 8004 15899 8007
rect 15887 7976 21772 8004
rect 15887 7973 15899 7976
rect 15841 7967 15899 7973
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7905 5779 7939
rect 8021 7939 8079 7945
rect 8021 7936 8033 7939
rect 5721 7899 5779 7905
rect 7208 7908 8033 7936
rect 7208 7880 7236 7908
rect 8021 7905 8033 7908
rect 8067 7905 8079 7939
rect 9582 7936 9588 7948
rect 8021 7899 8079 7905
rect 9508 7908 9588 7936
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4246 7868 4252 7880
rect 4203 7840 4252 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 5534 7828 5540 7880
rect 5592 7828 5598 7880
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 6822 7868 6828 7880
rect 6687 7840 6828 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7190 7828 7196 7880
rect 7248 7828 7254 7880
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7708 7840 7941 7868
rect 7708 7828 7714 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 9398 7868 9404 7880
rect 9355 7840 9404 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 9508 7877 9536 7908
rect 9582 7896 9588 7908
rect 9640 7936 9646 7948
rect 11057 7939 11115 7945
rect 11057 7936 11069 7939
rect 9640 7908 11069 7936
rect 9640 7896 9646 7908
rect 11057 7905 11069 7908
rect 11103 7905 11115 7939
rect 11057 7899 11115 7905
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11793 7939 11851 7945
rect 11793 7936 11805 7939
rect 11296 7908 11805 7936
rect 11296 7896 11302 7908
rect 11793 7905 11805 7908
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 13998 7936 14004 7948
rect 13320 7908 14004 7936
rect 13320 7896 13326 7908
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 14550 7896 14556 7948
rect 14608 7896 14614 7948
rect 16942 7896 16948 7948
rect 17000 7896 17006 7948
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 17644 7908 17693 7936
rect 17644 7896 17650 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7905 17831 7939
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 17773 7899 17831 7905
rect 18064 7908 18521 7936
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 4614 7800 4620 7812
rect 2746 7772 4620 7800
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 7837 7803 7895 7809
rect 7837 7769 7849 7803
rect 7883 7800 7895 7803
rect 8386 7800 8392 7812
rect 7883 7772 8392 7800
rect 7883 7769 7895 7772
rect 7837 7763 7895 7769
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 9416 7800 9444 7828
rect 9784 7800 9812 7831
rect 10318 7828 10324 7880
rect 10376 7828 10382 7880
rect 10410 7828 10416 7880
rect 10468 7828 10474 7880
rect 10594 7828 10600 7880
rect 10652 7828 10658 7880
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11388 7840 11989 7868
rect 11388 7828 11394 7840
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 9416 7772 9812 7800
rect 14752 7800 14780 7831
rect 14826 7828 14832 7880
rect 14884 7828 14890 7880
rect 15105 7871 15163 7877
rect 15105 7837 15117 7871
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15120 7800 15148 7831
rect 15286 7828 15292 7880
rect 15344 7828 15350 7880
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7868 15715 7871
rect 15703 7840 16436 7868
rect 15703 7837 15715 7840
rect 15657 7831 15715 7837
rect 15672 7800 15700 7831
rect 14752 7772 14964 7800
rect 15120 7772 15700 7800
rect 1762 7692 1768 7744
rect 1820 7692 1826 7744
rect 1854 7692 1860 7744
rect 1912 7692 1918 7744
rect 2590 7692 2596 7744
rect 2648 7692 2654 7744
rect 2682 7692 2688 7744
rect 2740 7692 2746 7744
rect 4525 7735 4583 7741
rect 4525 7701 4537 7735
rect 4571 7732 4583 7735
rect 5074 7732 5080 7744
rect 4571 7704 5080 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7732 5227 7735
rect 5350 7732 5356 7744
rect 5215 7704 5356 7732
rect 5215 7701 5227 7704
rect 5169 7695 5227 7701
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 6457 7735 6515 7741
rect 6457 7732 6469 7735
rect 5592 7704 6469 7732
rect 5592 7692 5598 7704
rect 6457 7701 6469 7704
rect 6503 7701 6515 7735
rect 6457 7695 6515 7701
rect 7374 7692 7380 7744
rect 7432 7692 7438 7744
rect 9950 7692 9956 7744
rect 10008 7692 10014 7744
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 12161 7735 12219 7741
rect 12161 7732 12173 7735
rect 10192 7704 12173 7732
rect 10192 7692 10198 7704
rect 12161 7701 12173 7704
rect 12207 7701 12219 7735
rect 12161 7695 12219 7701
rect 12986 7692 12992 7744
rect 13044 7692 13050 7744
rect 13078 7692 13084 7744
rect 13136 7692 13142 7744
rect 14936 7732 14964 7772
rect 15286 7732 15292 7744
rect 14936 7704 15292 7732
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 16408 7741 16436 7840
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17788 7868 17816 7899
rect 17862 7868 17868 7880
rect 17276 7840 17868 7868
rect 17276 7828 17282 7840
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 16761 7803 16819 7809
rect 16761 7769 16773 7803
rect 16807 7800 16819 7803
rect 17589 7803 17647 7809
rect 16807 7772 17540 7800
rect 16807 7769 16819 7772
rect 16761 7763 16819 7769
rect 16393 7735 16451 7741
rect 16393 7701 16405 7735
rect 16439 7701 16451 7735
rect 16393 7695 16451 7701
rect 16853 7735 16911 7741
rect 16853 7701 16865 7735
rect 16899 7732 16911 7735
rect 17221 7735 17279 7741
rect 17221 7732 17233 7735
rect 16899 7704 17233 7732
rect 16899 7701 16911 7704
rect 16853 7695 16911 7701
rect 17221 7701 17233 7704
rect 17267 7701 17279 7735
rect 17512 7732 17540 7772
rect 17589 7769 17601 7803
rect 17635 7800 17647 7803
rect 18064 7800 18092 7908
rect 18509 7905 18521 7908
rect 18555 7905 18567 7939
rect 18509 7899 18567 7905
rect 18969 7939 19027 7945
rect 18969 7905 18981 7939
rect 19015 7936 19027 7939
rect 19242 7936 19248 7948
rect 19015 7908 19248 7936
rect 19015 7905 19027 7908
rect 18969 7899 19027 7905
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19426 7868 19432 7880
rect 18923 7840 19432 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 17635 7772 18092 7800
rect 17635 7769 17647 7772
rect 17589 7763 17647 7769
rect 18138 7760 18144 7812
rect 18196 7800 18202 7812
rect 19812 7800 19840 7899
rect 21744 7877 21772 7976
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 18196 7772 19840 7800
rect 18196 7760 18202 7772
rect 19245 7735 19303 7741
rect 19245 7732 19257 7735
rect 17512 7704 19257 7732
rect 17221 7695 17279 7701
rect 19245 7701 19257 7704
rect 19291 7701 19303 7735
rect 19245 7695 19303 7701
rect 19610 7692 19616 7744
rect 19668 7692 19674 7744
rect 19705 7735 19763 7741
rect 19705 7701 19717 7735
rect 19751 7732 19763 7735
rect 19886 7732 19892 7744
rect 19751 7704 19892 7732
rect 19751 7701 19763 7704
rect 19705 7695 19763 7701
rect 19886 7692 19892 7704
rect 19944 7692 19950 7744
rect 21910 7692 21916 7744
rect 21968 7692 21974 7744
rect 1104 7642 22356 7664
rect 1104 7590 4266 7642
rect 4318 7590 4330 7642
rect 4382 7590 4394 7642
rect 4446 7590 4458 7642
rect 4510 7590 4522 7642
rect 4574 7590 9579 7642
rect 9631 7590 9643 7642
rect 9695 7590 9707 7642
rect 9759 7590 9771 7642
rect 9823 7590 9835 7642
rect 9887 7590 14892 7642
rect 14944 7590 14956 7642
rect 15008 7590 15020 7642
rect 15072 7590 15084 7642
rect 15136 7590 15148 7642
rect 15200 7590 20205 7642
rect 20257 7590 20269 7642
rect 20321 7590 20333 7642
rect 20385 7590 20397 7642
rect 20449 7590 20461 7642
rect 20513 7590 22356 7642
rect 1104 7568 22356 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 1596 7460 1624 7491
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2087 7531 2145 7537
rect 2087 7528 2099 7531
rect 1820 7500 2099 7528
rect 1820 7488 1826 7500
rect 2087 7497 2099 7500
rect 2133 7497 2145 7531
rect 2087 7491 2145 7497
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 2731 7531 2789 7537
rect 2731 7528 2743 7531
rect 2648 7500 2743 7528
rect 2648 7488 2654 7500
rect 2731 7497 2743 7500
rect 2777 7497 2789 7531
rect 2731 7491 2789 7497
rect 5350 7488 5356 7540
rect 5408 7488 5414 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 7190 7528 7196 7540
rect 5859 7500 7196 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 12986 7488 12992 7540
rect 13044 7528 13050 7540
rect 13173 7531 13231 7537
rect 13173 7528 13185 7531
rect 13044 7500 13185 7528
rect 13044 7488 13050 7500
rect 13173 7497 13185 7500
rect 13219 7497 13231 7531
rect 13173 7491 13231 7497
rect 18785 7531 18843 7537
rect 18785 7497 18797 7531
rect 18831 7528 18843 7531
rect 19610 7528 19616 7540
rect 18831 7500 19616 7528
rect 18831 7497 18843 7500
rect 18785 7491 18843 7497
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 2406 7460 2412 7472
rect 1596 7432 2412 7460
rect 2406 7420 2412 7432
rect 2464 7420 2470 7472
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 4433 7463 4491 7469
rect 4433 7460 4445 7463
rect 4212 7432 4445 7460
rect 4212 7420 4218 7432
rect 4433 7429 4445 7432
rect 4479 7429 4491 7463
rect 4433 7423 4491 7429
rect 5074 7420 5080 7472
rect 5132 7460 5138 7472
rect 5445 7463 5503 7469
rect 5445 7460 5457 7463
rect 5132 7432 5457 7460
rect 5132 7420 5138 7432
rect 5445 7429 5457 7432
rect 5491 7429 5503 7463
rect 5445 7423 5503 7429
rect 9950 7420 9956 7472
rect 10008 7420 10014 7472
rect 10134 7420 10140 7472
rect 10192 7420 10198 7472
rect 12713 7463 12771 7469
rect 12713 7429 12725 7463
rect 12759 7460 12771 7463
rect 13078 7460 13084 7472
rect 12759 7432 13084 7460
rect 12759 7429 12771 7432
rect 12713 7423 12771 7429
rect 13078 7420 13084 7432
rect 13136 7420 13142 7472
rect 18509 7463 18567 7469
rect 18509 7429 18521 7463
rect 18555 7460 18567 7463
rect 18966 7460 18972 7472
rect 18555 7432 18972 7460
rect 18555 7429 18567 7432
rect 18509 7423 18567 7429
rect 18966 7420 18972 7432
rect 19024 7420 19030 7472
rect 19334 7460 19340 7472
rect 19076 7432 19340 7460
rect 842 7352 848 7404
rect 900 7392 906 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 900 7364 1409 7392
rect 900 7352 906 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2158 7395 2216 7401
rect 2158 7392 2170 7395
rect 1912 7364 2170 7392
rect 1912 7352 1918 7364
rect 2158 7361 2170 7364
rect 2204 7361 2216 7395
rect 2158 7355 2216 7361
rect 2590 7352 2596 7404
rect 2648 7401 2654 7404
rect 2648 7395 2686 7401
rect 2674 7361 2686 7395
rect 2648 7355 2686 7361
rect 2648 7352 2654 7355
rect 3234 7352 3240 7404
rect 3292 7352 3298 7404
rect 4706 7392 4712 7404
rect 3620 7364 4712 7392
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 3620 7333 3648 7364
rect 4706 7352 4712 7364
rect 4764 7392 4770 7404
rect 4893 7395 4951 7401
rect 4893 7392 4905 7395
rect 4764 7364 4905 7392
rect 4764 7352 4770 7364
rect 4893 7361 4905 7364
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 7650 7352 7656 7404
rect 7708 7352 7714 7404
rect 12363 7395 12421 7401
rect 12363 7361 12375 7395
rect 12409 7392 12421 7395
rect 12409 7361 12434 7392
rect 12363 7355 12434 7361
rect 3145 7327 3203 7333
rect 3145 7324 3157 7327
rect 3108 7296 3157 7324
rect 3108 7284 3114 7296
rect 3145 7293 3157 7296
rect 3191 7293 3203 7327
rect 3145 7287 3203 7293
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4856 7296 4997 7324
rect 4856 7284 4862 7296
rect 4985 7293 4997 7296
rect 5031 7293 5043 7327
rect 4985 7287 5043 7293
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7324 5319 7327
rect 5994 7324 6000 7336
rect 5307 7296 6000 7324
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 12406 7324 12434 7355
rect 12526 7352 12532 7404
rect 12584 7392 12590 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12584 7364 13001 7392
rect 12584 7352 12590 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 14090 7352 14096 7404
rect 14148 7392 14154 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 14148 7364 14473 7392
rect 14148 7352 14154 7364
rect 14461 7361 14473 7364
rect 14507 7392 14519 7395
rect 14734 7392 14740 7404
rect 14507 7364 14740 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15194 7392 15200 7404
rect 15151 7364 15200 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 19076 7392 19104 7432
rect 19334 7420 19340 7432
rect 19392 7420 19398 7472
rect 20625 7463 20683 7469
rect 20625 7429 20637 7463
rect 20671 7460 20683 7463
rect 20671 7432 21312 7460
rect 20671 7429 20683 7432
rect 20625 7423 20683 7429
rect 21284 7401 21312 7432
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 18739 7364 19104 7392
rect 19168 7364 19625 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19168 7333 19196 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 21131 7395 21189 7401
rect 21131 7392 21143 7395
rect 20763 7364 21143 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 21131 7361 21143 7364
rect 21177 7361 21189 7395
rect 21131 7355 21189 7361
rect 21234 7395 21312 7401
rect 21234 7361 21246 7395
rect 21280 7361 21312 7395
rect 21234 7355 21312 7361
rect 21510 7395 21568 7401
rect 21510 7361 21522 7395
rect 21556 7392 21568 7395
rect 21818 7392 21824 7404
rect 21556 7364 21824 7392
rect 21556 7361 21568 7364
rect 21510 7355 21568 7361
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 12406 7296 12817 7324
rect 12406 7268 12434 7296
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 18969 7327 19027 7333
rect 18969 7293 18981 7327
rect 19015 7293 19027 7327
rect 18969 7287 19027 7293
rect 19153 7327 19211 7333
rect 19153 7293 19165 7327
rect 19199 7293 19211 7327
rect 19153 7287 19211 7293
rect 1854 7216 1860 7268
rect 1912 7216 1918 7268
rect 1946 7216 1952 7268
rect 2004 7256 2010 7268
rect 4154 7256 4160 7268
rect 2004 7228 4160 7256
rect 2004 7216 2010 7228
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 12342 7216 12348 7268
rect 12400 7228 12434 7268
rect 14645 7259 14703 7265
rect 12400 7216 12406 7228
rect 14645 7225 14657 7259
rect 14691 7256 14703 7259
rect 16758 7256 16764 7268
rect 14691 7228 16764 7256
rect 14691 7225 14703 7228
rect 14645 7219 14703 7225
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 18984 7256 19012 7287
rect 19242 7284 19248 7336
rect 19300 7284 19306 7336
rect 19521 7327 19579 7333
rect 19521 7293 19533 7327
rect 19567 7293 19579 7327
rect 19521 7287 19579 7293
rect 19426 7256 19432 7268
rect 18984 7228 19432 7256
rect 19426 7216 19432 7228
rect 19484 7256 19490 7268
rect 19536 7256 19564 7287
rect 19484 7228 19564 7256
rect 19628 7256 19656 7355
rect 19978 7284 19984 7336
rect 20036 7324 20042 7336
rect 20530 7324 20536 7336
rect 20036 7296 20536 7324
rect 20036 7284 20042 7296
rect 20530 7284 20536 7296
rect 20588 7324 20594 7336
rect 20809 7327 20867 7333
rect 20809 7324 20821 7327
rect 20588 7296 20821 7324
rect 20588 7284 20594 7296
rect 20809 7293 20821 7296
rect 20855 7293 20867 7327
rect 21284 7324 21312 7355
rect 21818 7352 21824 7364
rect 21876 7352 21882 7404
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 21284 7296 21864 7324
rect 20809 7287 20867 7293
rect 20254 7256 20260 7268
rect 19628 7228 20260 7256
rect 19484 7216 19490 7228
rect 20254 7216 20260 7228
rect 20312 7216 20318 7268
rect 21836 7265 21864 7296
rect 21821 7259 21879 7265
rect 21821 7225 21833 7259
rect 21867 7225 21879 7259
rect 21821 7219 21879 7225
rect 7834 7148 7840 7200
rect 7892 7148 7898 7200
rect 10318 7148 10324 7200
rect 10376 7148 10382 7200
rect 15289 7191 15347 7197
rect 15289 7157 15301 7191
rect 15335 7188 15347 7191
rect 15562 7188 15568 7200
rect 15335 7160 15568 7188
rect 15335 7157 15347 7160
rect 15289 7151 15347 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 18322 7148 18328 7200
rect 18380 7148 18386 7200
rect 20898 7148 20904 7200
rect 20956 7188 20962 7200
rect 21407 7191 21465 7197
rect 21407 7188 21419 7191
rect 20956 7160 21419 7188
rect 20956 7148 20962 7160
rect 21407 7157 21419 7160
rect 21453 7157 21465 7191
rect 21407 7151 21465 7157
rect 1104 7098 22356 7120
rect 1104 7046 3606 7098
rect 3658 7046 3670 7098
rect 3722 7046 3734 7098
rect 3786 7046 3798 7098
rect 3850 7046 3862 7098
rect 3914 7046 8919 7098
rect 8971 7046 8983 7098
rect 9035 7046 9047 7098
rect 9099 7046 9111 7098
rect 9163 7046 9175 7098
rect 9227 7046 14232 7098
rect 14284 7046 14296 7098
rect 14348 7046 14360 7098
rect 14412 7046 14424 7098
rect 14476 7046 14488 7098
rect 14540 7046 19545 7098
rect 19597 7046 19609 7098
rect 19661 7046 19673 7098
rect 19725 7046 19737 7098
rect 19789 7046 19801 7098
rect 19853 7046 22356 7098
rect 1104 7024 22356 7046
rect 6549 6987 6607 6993
rect 6549 6953 6561 6987
rect 6595 6984 6607 6987
rect 6822 6984 6828 6996
rect 6595 6956 6828 6984
rect 6595 6953 6607 6956
rect 6549 6947 6607 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 15565 6987 15623 6993
rect 15565 6984 15577 6987
rect 15252 6956 15577 6984
rect 15252 6944 15258 6956
rect 15565 6953 15577 6956
rect 15611 6953 15623 6987
rect 15565 6947 15623 6953
rect 19886 6944 19892 6996
rect 19944 6944 19950 6996
rect 17218 6876 17224 6928
rect 17276 6916 17282 6928
rect 20441 6919 20499 6925
rect 20441 6916 20453 6919
rect 17276 6888 18276 6916
rect 17276 6876 17282 6888
rect 5258 6808 5264 6860
rect 5316 6808 5322 6860
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6546 6848 6552 6860
rect 6052 6820 6552 6848
rect 6052 6808 6058 6820
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 12618 6808 12624 6860
rect 12676 6808 12682 6860
rect 13078 6808 13084 6860
rect 13136 6808 13142 6860
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 15838 6848 15844 6860
rect 14700 6820 15844 6848
rect 14700 6808 14706 6820
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16114 6808 16120 6860
rect 16172 6848 16178 6860
rect 16942 6848 16948 6860
rect 16172 6820 16948 6848
rect 16172 6808 16178 6820
rect 16942 6808 16948 6820
rect 17000 6848 17006 6860
rect 18248 6857 18276 6888
rect 20088 6888 20453 6916
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 17000 6820 17417 6848
rect 17000 6808 17006 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 18233 6851 18291 6857
rect 18233 6817 18245 6851
rect 18279 6817 18291 6851
rect 18233 6811 18291 6817
rect 18322 6808 18328 6860
rect 18380 6848 18386 6860
rect 19058 6848 19064 6860
rect 18380 6820 19064 6848
rect 18380 6808 18386 6820
rect 19058 6808 19064 6820
rect 19116 6848 19122 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 19116 6820 19257 6848
rect 19116 6808 19122 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 5276 6780 5304 6808
rect 5442 6780 5448 6792
rect 5276 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6780 5506 6792
rect 5500 6752 6408 6780
rect 5500 6740 5506 6752
rect 5074 6672 5080 6724
rect 5132 6672 5138 6724
rect 5258 6672 5264 6724
rect 5316 6712 5322 6724
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 5316 6684 6193 6712
rect 5316 6672 5322 6684
rect 6181 6681 6193 6684
rect 6227 6681 6239 6715
rect 6380 6712 6408 6752
rect 6822 6740 6828 6792
rect 6880 6740 6886 6792
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6780 13047 6783
rect 13906 6780 13912 6792
rect 13035 6752 13912 6780
rect 13035 6749 13047 6752
rect 12989 6743 13047 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14660 6712 14688 6808
rect 20088 6792 20116 6888
rect 20441 6885 20453 6888
rect 20487 6885 20499 6919
rect 20441 6879 20499 6885
rect 20714 6876 20720 6928
rect 20772 6916 20778 6928
rect 20772 6888 21036 6916
rect 20772 6876 20778 6888
rect 20898 6808 20904 6860
rect 20956 6808 20962 6860
rect 21008 6857 21036 6888
rect 20993 6851 21051 6857
rect 20993 6817 21005 6851
rect 21039 6817 21051 6851
rect 20993 6811 21051 6817
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6780 18199 6783
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 18187 6752 18521 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 18509 6749 18521 6752
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 20070 6780 20076 6792
rect 19484 6752 20076 6780
rect 19484 6740 19490 6752
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 20254 6740 20260 6792
rect 20312 6780 20318 6792
rect 20530 6780 20536 6792
rect 20312 6752 20536 6780
rect 20312 6740 20318 6752
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 6380 6684 14688 6712
rect 15933 6715 15991 6721
rect 6181 6675 6239 6681
rect 15933 6681 15945 6715
rect 15979 6712 15991 6715
rect 16574 6712 16580 6724
rect 15979 6684 16580 6712
rect 15979 6681 15991 6684
rect 15933 6675 15991 6681
rect 16574 6672 16580 6684
rect 16632 6672 16638 6724
rect 17221 6715 17279 6721
rect 17221 6681 17233 6715
rect 17267 6712 17279 6715
rect 18230 6712 18236 6724
rect 17267 6684 18236 6712
rect 17267 6681 17279 6684
rect 17221 6675 17279 6681
rect 18230 6672 18236 6684
rect 18288 6672 18294 6724
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 5534 6644 5540 6656
rect 3384 6616 5540 6644
rect 3384 6604 3390 6616
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 6086 6604 6092 6656
rect 6144 6604 6150 6656
rect 8570 6604 8576 6656
rect 8628 6604 8634 6656
rect 16025 6647 16083 6653
rect 16025 6613 16037 6647
rect 16071 6644 16083 6647
rect 16666 6644 16672 6656
rect 16071 6616 16672 6644
rect 16071 6613 16083 6616
rect 16025 6607 16083 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 17126 6644 17132 6656
rect 16899 6616 17132 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 17313 6647 17371 6653
rect 17313 6613 17325 6647
rect 17359 6644 17371 6647
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17359 6616 17693 6644
rect 17359 6613 17371 6616
rect 17313 6607 17371 6613
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17681 6607 17739 6613
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6644 18107 6647
rect 18414 6644 18420 6656
rect 18095 6616 18420 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 18782 6604 18788 6656
rect 18840 6644 18846 6656
rect 19705 6647 19763 6653
rect 19705 6644 19717 6647
rect 18840 6616 19717 6644
rect 18840 6604 18846 6616
rect 19705 6613 19717 6616
rect 19751 6613 19763 6647
rect 19705 6607 19763 6613
rect 20809 6647 20867 6653
rect 20809 6613 20821 6647
rect 20855 6644 20867 6647
rect 21818 6644 21824 6656
rect 20855 6616 21824 6644
rect 20855 6613 20867 6616
rect 20809 6607 20867 6613
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 1104 6554 22356 6576
rect 1104 6502 4266 6554
rect 4318 6502 4330 6554
rect 4382 6502 4394 6554
rect 4446 6502 4458 6554
rect 4510 6502 4522 6554
rect 4574 6502 9579 6554
rect 9631 6502 9643 6554
rect 9695 6502 9707 6554
rect 9759 6502 9771 6554
rect 9823 6502 9835 6554
rect 9887 6502 14892 6554
rect 14944 6502 14956 6554
rect 15008 6502 15020 6554
rect 15072 6502 15084 6554
rect 15136 6502 15148 6554
rect 15200 6502 20205 6554
rect 20257 6502 20269 6554
rect 20321 6502 20333 6554
rect 20385 6502 20397 6554
rect 20449 6502 20461 6554
rect 20513 6502 22356 6554
rect 1104 6480 22356 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 2590 6440 2596 6452
rect 1627 6412 2596 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 4798 6440 4804 6452
rect 4479 6412 4804 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 5258 6400 5264 6452
rect 5316 6400 5322 6452
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 6144 6412 6377 6440
rect 6144 6400 6150 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6822 6400 6828 6452
rect 6880 6400 6886 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7708 6412 8033 6440
rect 7708 6400 7714 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 8021 6403 8079 6409
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8444 6412 8861 6440
rect 8444 6400 8450 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 9355 6412 9689 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 9677 6403 9735 6409
rect 16666 6400 16672 6452
rect 16724 6400 16730 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19889 6443 19947 6449
rect 19889 6440 19901 6443
rect 19392 6412 19901 6440
rect 19392 6400 19398 6412
rect 19889 6409 19901 6412
rect 19935 6409 19947 6443
rect 19889 6403 19947 6409
rect 4249 6375 4307 6381
rect 4249 6341 4261 6375
rect 4295 6372 4307 6375
rect 4982 6372 4988 6384
rect 4295 6344 4988 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 4982 6332 4988 6344
rect 5040 6332 5046 6384
rect 5442 6332 5448 6384
rect 5500 6332 5506 6384
rect 14642 6332 14648 6384
rect 14700 6332 14706 6384
rect 14737 6375 14795 6381
rect 14737 6341 14749 6375
rect 14783 6372 14795 6375
rect 16114 6372 16120 6384
rect 14783 6344 16120 6372
rect 14783 6341 14795 6344
rect 14737 6335 14795 6341
rect 16114 6332 16120 6344
rect 16172 6332 16178 6384
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 3510 6264 3516 6316
rect 3568 6304 3574 6316
rect 3732 6307 3790 6313
rect 3732 6304 3744 6307
rect 3568 6276 3744 6304
rect 3568 6264 3574 6276
rect 3732 6273 3744 6276
rect 3778 6273 3790 6307
rect 3732 6267 3790 6273
rect 3970 6264 3976 6316
rect 4028 6304 4034 6316
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 4028 6276 4077 6304
rect 4028 6264 4034 6276
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 4212 6276 4905 6304
rect 4212 6264 4218 6276
rect 4893 6273 4905 6276
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6144 6276 6745 6304
rect 6144 6264 6150 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 7650 6264 7656 6316
rect 7708 6264 7714 6316
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9490 6304 9496 6316
rect 9263 6276 9496 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 9766 6264 9772 6316
rect 9824 6304 9830 6316
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9824 6276 10057 6304
rect 9824 6264 9830 6276
rect 10045 6273 10057 6276
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10183 6276 10517 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 12066 6264 12072 6316
rect 12124 6304 12130 6316
rect 12342 6304 12348 6316
rect 12124 6276 12348 6304
rect 12124 6264 12130 6276
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12728 6276 13001 6304
rect 4706 6196 4712 6248
rect 4764 6196 4770 6248
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 4816 6112 4844 6199
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5408 6208 5733 6236
rect 5408 6196 5414 6208
rect 5721 6205 5733 6208
rect 5767 6236 5779 6239
rect 7006 6236 7012 6248
rect 5767 6208 7012 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 4890 6128 4896 6180
rect 4948 6168 4954 6180
rect 5368 6168 5396 6196
rect 4948 6140 5396 6168
rect 4948 6128 4954 6140
rect 6546 6128 6552 6180
rect 6604 6168 6610 6180
rect 7484 6168 7512 6199
rect 7558 6196 7564 6248
rect 7616 6196 7622 6248
rect 9398 6196 9404 6248
rect 9456 6196 9462 6248
rect 10226 6196 10232 6248
rect 10284 6196 10290 6248
rect 12728 6245 12756 6276
rect 12989 6273 13001 6276
rect 13035 6304 13047 6307
rect 13078 6304 13084 6316
rect 13035 6276 13084 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6304 13507 6307
rect 13814 6304 13820 6316
rect 13495 6276 13820 6304
rect 13495 6273 13507 6276
rect 13449 6267 13507 6273
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 17034 6264 17040 6316
rect 17092 6264 17098 6316
rect 18782 6264 18788 6316
rect 18840 6264 18846 6316
rect 20070 6264 20076 6316
rect 20128 6264 20134 6316
rect 21174 6264 21180 6316
rect 21232 6304 21238 6316
rect 21361 6307 21419 6313
rect 21361 6304 21373 6307
rect 21232 6276 21373 6304
rect 21232 6264 21238 6276
rect 21361 6273 21373 6276
rect 21407 6273 21419 6307
rect 21361 6267 21419 6273
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 12437 6239 12495 6245
rect 11931 6208 12204 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 9416 6168 9444 6196
rect 6604 6140 9444 6168
rect 6604 6128 6610 6140
rect 12066 6128 12072 6180
rect 12124 6128 12130 6180
rect 12176 6168 12204 6208
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12713 6239 12771 6245
rect 12483 6208 12517 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12713 6205 12725 6239
rect 12759 6205 12771 6239
rect 12713 6199 12771 6205
rect 12805 6239 12863 6245
rect 12805 6205 12817 6239
rect 12851 6236 12863 6239
rect 13541 6239 13599 6245
rect 13541 6236 13553 6239
rect 12851 6208 13553 6236
rect 12851 6205 12863 6208
rect 12805 6199 12863 6205
rect 13541 6205 13553 6208
rect 13587 6236 13599 6239
rect 13906 6236 13912 6248
rect 13587 6208 13912 6236
rect 13587 6205 13599 6208
rect 13541 6199 13599 6205
rect 12452 6168 12480 6199
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 14550 6196 14556 6248
rect 14608 6196 14614 6248
rect 16485 6239 16543 6245
rect 16485 6205 16497 6239
rect 16531 6236 16543 6239
rect 17129 6239 17187 6245
rect 17129 6236 17141 6239
rect 16531 6208 17141 6236
rect 16531 6205 16543 6208
rect 16485 6199 16543 6205
rect 17129 6205 17141 6208
rect 17175 6205 17187 6239
rect 17129 6199 17187 6205
rect 17218 6196 17224 6248
rect 17276 6196 17282 6248
rect 18414 6196 18420 6248
rect 18472 6196 18478 6248
rect 18874 6196 18880 6248
rect 18932 6196 18938 6248
rect 20257 6239 20315 6245
rect 20257 6205 20269 6239
rect 20303 6236 20315 6239
rect 20530 6236 20536 6248
rect 20303 6208 20536 6236
rect 20303 6205 20315 6208
rect 20257 6199 20315 6205
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 12526 6168 12532 6180
rect 12176 6140 12532 6168
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 14090 6128 14096 6180
rect 14148 6168 14154 6180
rect 14185 6171 14243 6177
rect 14185 6168 14197 6171
rect 14148 6140 14197 6168
rect 14148 6128 14154 6140
rect 14185 6137 14197 6140
rect 14231 6137 14243 6171
rect 18782 6168 18788 6180
rect 14185 6131 14243 6137
rect 14844 6140 18788 6168
rect 3835 6103 3893 6109
rect 3835 6069 3847 6103
rect 3881 6100 3893 6103
rect 4062 6100 4068 6112
rect 3881 6072 4068 6100
rect 3881 6069 3893 6072
rect 3835 6063 3893 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4798 6060 4804 6112
rect 4856 6060 4862 6112
rect 8110 6060 8116 6112
rect 8168 6060 8174 6112
rect 11701 6103 11759 6109
rect 11701 6069 11713 6103
rect 11747 6100 11759 6103
rect 12986 6100 12992 6112
rect 11747 6072 12992 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13170 6060 13176 6112
rect 13228 6060 13234 6112
rect 13817 6103 13875 6109
rect 13817 6069 13829 6103
rect 13863 6100 13875 6103
rect 14844 6100 14872 6140
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 21542 6128 21548 6180
rect 21600 6128 21606 6180
rect 13863 6072 14872 6100
rect 13863 6069 13875 6072
rect 13817 6063 13875 6069
rect 14918 6060 14924 6112
rect 14976 6060 14982 6112
rect 1104 6010 22356 6032
rect 1104 5958 3606 6010
rect 3658 5958 3670 6010
rect 3722 5958 3734 6010
rect 3786 5958 3798 6010
rect 3850 5958 3862 6010
rect 3914 5958 8919 6010
rect 8971 5958 8983 6010
rect 9035 5958 9047 6010
rect 9099 5958 9111 6010
rect 9163 5958 9175 6010
rect 9227 5958 14232 6010
rect 14284 5958 14296 6010
rect 14348 5958 14360 6010
rect 14412 5958 14424 6010
rect 14476 5958 14488 6010
rect 14540 5958 19545 6010
rect 19597 5958 19609 6010
rect 19661 5958 19673 6010
rect 19725 5958 19737 6010
rect 19789 5958 19801 6010
rect 19853 5958 22356 6010
rect 1104 5936 22356 5958
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 3970 5896 3976 5908
rect 3283 5868 3976 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 6086 5856 6092 5908
rect 6144 5856 6150 5908
rect 7558 5856 7564 5908
rect 7616 5856 7622 5908
rect 8110 5856 8116 5908
rect 8168 5856 8174 5908
rect 9766 5856 9772 5908
rect 9824 5856 9830 5908
rect 10686 5856 10692 5908
rect 10744 5856 10750 5908
rect 11885 5899 11943 5905
rect 11885 5865 11897 5899
rect 11931 5896 11943 5899
rect 12526 5896 12532 5908
rect 11931 5868 12532 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 12526 5856 12532 5868
rect 12584 5856 12590 5908
rect 14461 5899 14519 5905
rect 14461 5865 14473 5899
rect 14507 5896 14519 5899
rect 14642 5896 14648 5908
rect 14507 5868 14648 5896
rect 14507 5865 14519 5868
rect 14461 5859 14519 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 21818 5856 21824 5908
rect 21876 5856 21882 5908
rect 3605 5831 3663 5837
rect 3605 5797 3617 5831
rect 3651 5828 3663 5831
rect 4525 5831 4583 5837
rect 4525 5828 4537 5831
rect 3651 5800 4537 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 4525 5797 4537 5800
rect 4571 5797 4583 5831
rect 8128 5828 8156 5856
rect 10226 5828 10232 5840
rect 4525 5791 4583 5797
rect 8036 5800 8156 5828
rect 8220 5800 10232 5828
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 4246 5760 4252 5772
rect 3927 5732 4252 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 3326 5692 3332 5704
rect 1719 5664 3332 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3970 5692 3976 5704
rect 3467 5664 3976 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4540 5692 4568 5791
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5760 5227 5763
rect 5442 5760 5448 5772
rect 5215 5732 5448 5760
rect 5215 5729 5227 5732
rect 5169 5723 5227 5729
rect 4614 5692 4620 5704
rect 4540 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5692 4678 5704
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4672 5664 4813 5692
rect 4672 5652 4678 5664
rect 4801 5661 4813 5664
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 3988 5624 4016 5652
rect 4908 5624 4936 5723
rect 5442 5720 5448 5732
rect 5500 5760 5506 5772
rect 8036 5769 8064 5800
rect 8220 5769 8248 5800
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 13998 5788 14004 5840
rect 14056 5828 14062 5840
rect 14056 5800 15056 5828
rect 14056 5788 14062 5800
rect 5629 5763 5687 5769
rect 5629 5760 5641 5763
rect 5500 5732 5641 5760
rect 5500 5720 5506 5732
rect 5629 5729 5641 5732
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 5718 5652 5724 5704
rect 5776 5652 5782 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7190 5692 7196 5704
rect 7064 5664 7196 5692
rect 7064 5652 7070 5664
rect 7190 5652 7196 5664
rect 7248 5692 7254 5704
rect 8220 5692 8248 5723
rect 10042 5720 10048 5772
rect 10100 5720 10106 5772
rect 10318 5760 10324 5772
rect 10152 5732 10324 5760
rect 10152 5701 10180 5732
rect 10318 5720 10324 5732
rect 10376 5760 10382 5772
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 10376 5732 10425 5760
rect 10376 5720 10382 5732
rect 10413 5729 10425 5732
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 11790 5720 11796 5772
rect 11848 5760 11854 5772
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 11848 5732 12449 5760
rect 11848 5720 11854 5732
rect 12437 5729 12449 5732
rect 12483 5729 12495 5763
rect 12437 5723 12495 5729
rect 14918 5720 14924 5772
rect 14976 5720 14982 5772
rect 15028 5769 15056 5800
rect 19058 5788 19064 5840
rect 19116 5788 19122 5840
rect 15013 5763 15071 5769
rect 15013 5729 15025 5763
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 7248 5664 8248 5692
rect 10137 5695 10195 5701
rect 7248 5652 7254 5664
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10505 5695 10563 5701
rect 10505 5661 10517 5695
rect 10551 5661 10563 5695
rect 10505 5655 10563 5661
rect 11676 5695 11734 5701
rect 11676 5661 11688 5695
rect 11722 5692 11734 5695
rect 12066 5692 12072 5704
rect 11722 5664 12072 5692
rect 11722 5661 11734 5664
rect 11676 5655 11734 5661
rect 3988 5596 4936 5624
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10520 5624 10548 5655
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12830 5695 12888 5701
rect 12830 5692 12842 5695
rect 12544 5664 12842 5692
rect 12544 5636 12572 5664
rect 12830 5661 12842 5664
rect 12876 5661 12888 5695
rect 12830 5655 12888 5661
rect 12986 5652 12992 5704
rect 13044 5652 13050 5704
rect 13170 5652 13176 5704
rect 13228 5652 13234 5704
rect 18874 5652 18880 5704
rect 18932 5652 18938 5704
rect 22002 5652 22008 5704
rect 22060 5652 22066 5704
rect 10100 5596 10548 5624
rect 12253 5627 12311 5633
rect 10100 5584 10106 5596
rect 12253 5593 12265 5627
rect 12299 5624 12311 5627
rect 12526 5624 12532 5636
rect 12299 5596 12532 5624
rect 12299 5593 12311 5596
rect 12253 5587 12311 5593
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 1486 5516 1492 5568
rect 1544 5516 1550 5568
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4157 5559 4215 5565
rect 4157 5556 4169 5559
rect 4120 5528 4169 5556
rect 4120 5516 4126 5528
rect 4157 5525 4169 5528
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 7558 5556 7564 5568
rect 4304 5528 7564 5556
rect 4304 5516 4310 5528
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 7926 5516 7932 5568
rect 7984 5516 7990 5568
rect 11790 5565 11796 5568
rect 11747 5559 11796 5565
rect 11747 5525 11759 5559
rect 11793 5525 11796 5559
rect 11747 5519 11796 5525
rect 11790 5516 11796 5519
rect 11848 5516 11854 5568
rect 12345 5559 12403 5565
rect 12345 5525 12357 5559
rect 12391 5556 12403 5559
rect 12759 5559 12817 5565
rect 12759 5556 12771 5559
rect 12391 5528 12771 5556
rect 12391 5525 12403 5528
rect 12345 5519 12403 5525
rect 12759 5525 12771 5528
rect 12805 5525 12817 5559
rect 12759 5519 12817 5525
rect 13357 5559 13415 5565
rect 13357 5525 13369 5559
rect 13403 5556 13415 5559
rect 13814 5556 13820 5568
rect 13403 5528 13820 5556
rect 13403 5525 13415 5528
rect 13357 5519 13415 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14734 5516 14740 5568
rect 14792 5556 14798 5568
rect 14829 5559 14887 5565
rect 14829 5556 14841 5559
rect 14792 5528 14841 5556
rect 14792 5516 14798 5528
rect 14829 5525 14841 5528
rect 14875 5525 14887 5559
rect 14829 5519 14887 5525
rect 18690 5516 18696 5568
rect 18748 5516 18754 5568
rect 1104 5466 22356 5488
rect 1104 5414 4266 5466
rect 4318 5414 4330 5466
rect 4382 5414 4394 5466
rect 4446 5414 4458 5466
rect 4510 5414 4522 5466
rect 4574 5414 9579 5466
rect 9631 5414 9643 5466
rect 9695 5414 9707 5466
rect 9759 5414 9771 5466
rect 9823 5414 9835 5466
rect 9887 5414 14892 5466
rect 14944 5414 14956 5466
rect 15008 5414 15020 5466
rect 15072 5414 15084 5466
rect 15136 5414 15148 5466
rect 15200 5414 20205 5466
rect 20257 5414 20269 5466
rect 20321 5414 20333 5466
rect 20385 5414 20397 5466
rect 20449 5414 20461 5466
rect 20513 5414 22356 5466
rect 1104 5392 22356 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 3510 5352 3516 5364
rect 1627 5324 3516 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 3510 5312 3516 5324
rect 3568 5352 3574 5364
rect 4062 5352 4068 5364
rect 3568 5324 4068 5352
rect 3568 5312 3574 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 4212 5324 4261 5352
rect 4212 5312 4218 5324
rect 4249 5321 4261 5324
rect 4295 5321 4307 5355
rect 4249 5315 4307 5321
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 4798 5352 4804 5364
rect 4755 5324 4804 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 11977 5355 12035 5361
rect 11977 5352 11989 5355
rect 11848 5324 11989 5352
rect 11848 5312 11854 5324
rect 11977 5321 11989 5324
rect 12023 5321 12035 5355
rect 11977 5315 12035 5321
rect 12342 5312 12348 5364
rect 12400 5352 12406 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 12400 5324 12449 5352
rect 12400 5312 12406 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 12437 5315 12495 5321
rect 18230 5312 18236 5364
rect 18288 5312 18294 5364
rect 21266 5312 21272 5364
rect 21324 5352 21330 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 21324 5324 21833 5352
rect 21324 5312 21330 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 4614 5284 4620 5296
rect 4387 5256 4620 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 4356 5216 4384 5247
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 4982 5244 4988 5296
rect 5040 5244 5046 5296
rect 7009 5287 7067 5293
rect 7009 5253 7021 5287
rect 7055 5284 7067 5287
rect 8389 5287 8447 5293
rect 8389 5284 8401 5287
rect 7055 5256 8401 5284
rect 7055 5253 7067 5256
rect 7009 5247 7067 5253
rect 8389 5253 8401 5256
rect 8435 5253 8447 5287
rect 8389 5247 8447 5253
rect 9769 5287 9827 5293
rect 9769 5253 9781 5287
rect 9815 5284 9827 5287
rect 10686 5284 10692 5296
rect 9815 5256 10692 5284
rect 9815 5253 9827 5256
rect 9769 5247 9827 5253
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 17218 5244 17224 5296
rect 17276 5284 17282 5296
rect 17276 5256 18828 5284
rect 17276 5244 17282 5256
rect 1397 5179 1455 5185
rect 3896 5188 4384 5216
rect 4525 5219 4583 5225
rect 3896 5157 3924 5188
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5117 3939 5151
rect 3881 5111 3939 5117
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 4065 5151 4123 5157
rect 4065 5148 4077 5151
rect 4028 5120 4077 5148
rect 4028 5108 4034 5120
rect 4065 5117 4077 5120
rect 4111 5148 4123 5151
rect 4540 5148 4568 5179
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7607 5188 8248 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 4111 5120 4568 5148
rect 5537 5151 5595 5157
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 5718 5148 5724 5160
rect 5583 5120 5724 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 5718 5108 5724 5120
rect 5776 5148 5782 5160
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 5776 5120 7205 5148
rect 5776 5108 5782 5120
rect 7193 5117 7205 5120
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 7469 5151 7527 5157
rect 7469 5148 7481 5151
rect 7340 5120 7481 5148
rect 7340 5108 7346 5120
rect 7469 5117 7481 5120
rect 7515 5117 7527 5151
rect 7469 5111 7527 5117
rect 7484 5080 7512 5111
rect 7926 5108 7932 5160
rect 7984 5108 7990 5160
rect 8220 5157 8248 5188
rect 9582 5176 9588 5228
rect 9640 5176 9646 5228
rect 12066 5176 12072 5228
rect 12124 5176 12130 5228
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 14148 5188 14381 5216
rect 14148 5176 14154 5188
rect 14369 5185 14381 5188
rect 14415 5216 14427 5219
rect 15102 5216 15108 5228
rect 14415 5188 15108 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5216 16911 5219
rect 16899 5188 17448 5216
rect 16899 5185 16911 5188
rect 16853 5179 16911 5185
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 8251 5120 9965 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 11885 5151 11943 5157
rect 11885 5117 11897 5151
rect 11931 5148 11943 5151
rect 11974 5148 11980 5160
rect 11931 5120 11980 5148
rect 11931 5117 11943 5120
rect 11885 5111 11943 5117
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 13722 5108 13728 5160
rect 13780 5148 13786 5160
rect 13909 5151 13967 5157
rect 13909 5148 13921 5151
rect 13780 5120 13921 5148
rect 13780 5108 13786 5120
rect 13909 5117 13921 5120
rect 13955 5117 13967 5151
rect 13909 5111 13967 5117
rect 14461 5151 14519 5157
rect 14461 5117 14473 5151
rect 14507 5148 14519 5151
rect 14642 5148 14648 5160
rect 14507 5120 14648 5148
rect 14507 5117 14519 5120
rect 14461 5111 14519 5117
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 16666 5108 16672 5160
rect 16724 5148 16730 5160
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 16724 5120 16773 5148
rect 16724 5108 16730 5120
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 17034 5108 17040 5160
rect 17092 5148 17098 5160
rect 17221 5151 17279 5157
rect 17221 5148 17233 5151
rect 17092 5120 17233 5148
rect 17092 5108 17098 5120
rect 17221 5117 17233 5120
rect 17267 5117 17279 5151
rect 17221 5111 17279 5117
rect 17420 5089 17448 5188
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 17736 5188 18613 5216
rect 17736 5176 17742 5188
rect 18601 5185 18613 5188
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 17862 5108 17868 5160
rect 17920 5108 17926 5160
rect 18800 5157 18828 5256
rect 19150 5176 19156 5228
rect 19208 5216 19214 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 19208 5188 19441 5216
rect 19208 5176 19214 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 22002 5176 22008 5228
rect 22060 5176 22066 5228
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18785 5151 18843 5157
rect 18785 5117 18797 5151
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 8021 5083 8079 5089
rect 8021 5080 8033 5083
rect 7484 5052 8033 5080
rect 8021 5049 8033 5052
rect 8067 5049 8079 5083
rect 8021 5043 8079 5049
rect 17405 5083 17463 5089
rect 17405 5049 17417 5083
rect 17451 5049 17463 5083
rect 18708 5080 18736 5111
rect 18874 5108 18880 5160
rect 18932 5148 18938 5160
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 18932 5120 19073 5148
rect 18932 5108 18938 5120
rect 19061 5117 19073 5120
rect 19107 5117 19119 5151
rect 19061 5111 19119 5117
rect 19334 5108 19340 5160
rect 19392 5108 19398 5160
rect 19242 5080 19248 5092
rect 18708 5052 19248 5080
rect 17405 5043 17463 5049
rect 19242 5040 19248 5052
rect 19300 5040 19306 5092
rect 1104 4922 22356 4944
rect 1104 4870 3606 4922
rect 3658 4870 3670 4922
rect 3722 4870 3734 4922
rect 3786 4870 3798 4922
rect 3850 4870 3862 4922
rect 3914 4870 8919 4922
rect 8971 4870 8983 4922
rect 9035 4870 9047 4922
rect 9099 4870 9111 4922
rect 9163 4870 9175 4922
rect 9227 4870 14232 4922
rect 14284 4870 14296 4922
rect 14348 4870 14360 4922
rect 14412 4870 14424 4922
rect 14476 4870 14488 4922
rect 14540 4870 19545 4922
rect 19597 4870 19609 4922
rect 19661 4870 19673 4922
rect 19725 4870 19737 4922
rect 19789 4870 19801 4922
rect 19853 4870 22356 4922
rect 1104 4848 22356 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 5074 4808 5080 4820
rect 1627 4780 5080 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4808 9091 4811
rect 9582 4808 9588 4820
rect 9079 4780 9588 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 10100 4780 10333 4808
rect 10100 4768 10106 4780
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 10321 4771 10379 4777
rect 13906 4768 13912 4820
rect 13964 4768 13970 4820
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 14792 4780 15117 4808
rect 14792 4768 14798 4780
rect 15105 4777 15117 4780
rect 15151 4777 15163 4811
rect 15105 4771 15163 4777
rect 17678 4768 17684 4820
rect 17736 4768 17742 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 18969 4811 19027 4817
rect 18969 4808 18981 4811
rect 17920 4780 18981 4808
rect 17920 4768 17926 4780
rect 18969 4777 18981 4780
rect 19015 4777 19027 4811
rect 18969 4771 19027 4777
rect 19242 4768 19248 4820
rect 19300 4768 19306 4820
rect 9490 4700 9496 4752
rect 9548 4700 9554 4752
rect 17313 4743 17371 4749
rect 17313 4740 17325 4743
rect 9968 4712 10916 4740
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 4764 4644 5825 4672
rect 4764 4632 4770 4644
rect 5813 4641 5825 4644
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 5626 4564 5632 4616
rect 5684 4564 5690 4616
rect 5828 4536 5856 4635
rect 7006 4632 7012 4684
rect 7064 4632 7070 4684
rect 9398 4632 9404 4684
rect 9456 4672 9462 4684
rect 9968 4672 9996 4712
rect 9456 4644 9996 4672
rect 10137 4675 10195 4681
rect 9456 4632 9462 4644
rect 10137 4641 10149 4675
rect 10183 4672 10195 4675
rect 10226 4672 10232 4684
rect 10183 4644 10232 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10778 4672 10784 4684
rect 10336 4644 10784 4672
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6972 4576 7205 4604
rect 6972 4564 6978 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 10336 4604 10364 4644
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 9263 4576 10364 4604
rect 10689 4607 10747 4613
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 10888 4604 10916 4712
rect 15396 4712 17325 4740
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4672 14519 4675
rect 14642 4672 14648 4684
rect 14507 4644 14648 4672
rect 14507 4641 14519 4644
rect 14461 4635 14519 4641
rect 14642 4632 14648 4644
rect 14700 4672 14706 4684
rect 15396 4672 15424 4712
rect 17313 4709 17325 4712
rect 17359 4709 17371 4743
rect 17313 4703 17371 4709
rect 14700 4644 15424 4672
rect 15565 4675 15623 4681
rect 14700 4632 14706 4644
rect 15565 4641 15577 4675
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 16853 4675 16911 4681
rect 16853 4641 16865 4675
rect 16899 4672 16911 4675
rect 17880 4672 17908 4768
rect 18049 4743 18107 4749
rect 18049 4709 18061 4743
rect 18095 4740 18107 4743
rect 18141 4743 18199 4749
rect 18141 4740 18153 4743
rect 18095 4712 18153 4740
rect 18095 4709 18107 4712
rect 18049 4703 18107 4709
rect 18141 4709 18153 4712
rect 18187 4740 18199 4743
rect 19150 4740 19156 4752
rect 18187 4712 19156 4740
rect 18187 4709 18199 4712
rect 18141 4703 18199 4709
rect 19150 4700 19156 4712
rect 19208 4700 19214 4752
rect 16899 4644 17908 4672
rect 18325 4675 18383 4681
rect 16899 4641 16911 4644
rect 16853 4635 16911 4641
rect 18325 4641 18337 4675
rect 18371 4672 18383 4675
rect 19334 4672 19340 4684
rect 18371 4644 19340 4672
rect 18371 4641 18383 4644
rect 18325 4635 18383 4641
rect 10735 4576 10916 4604
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 13722 4564 13728 4616
rect 13780 4564 13786 4616
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 14936 4576 15485 4604
rect 7742 4536 7748 4548
rect 5828 4508 7748 4536
rect 7742 4496 7748 4508
rect 7800 4496 7806 4548
rect 9861 4539 9919 4545
rect 9861 4505 9873 4539
rect 9907 4536 9919 4539
rect 10134 4536 10140 4548
rect 9907 4508 10140 4536
rect 9907 4505 9919 4508
rect 9861 4499 9919 4505
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 13538 4496 13544 4548
rect 13596 4496 13602 4548
rect 7377 4471 7435 4477
rect 7377 4437 7389 4471
rect 7423 4468 7435 4471
rect 7466 4468 7472 4480
rect 7423 4440 7472 4468
rect 7423 4437 7435 4440
rect 7377 4431 7435 4437
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 9950 4428 9956 4480
rect 10008 4428 10014 4480
rect 14936 4477 14964 4576
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 15102 4496 15108 4548
rect 15160 4536 15166 4548
rect 15580 4536 15608 4635
rect 15838 4564 15844 4616
rect 15896 4564 15902 4616
rect 16666 4564 16672 4616
rect 16724 4564 16730 4616
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4604 17923 4607
rect 18340 4604 18368 4635
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 20625 4675 20683 4681
rect 20625 4641 20637 4675
rect 20671 4672 20683 4675
rect 20714 4672 20720 4684
rect 20671 4644 20720 4672
rect 20671 4641 20683 4644
rect 20625 4635 20683 4641
rect 20714 4632 20720 4644
rect 20772 4632 20778 4684
rect 17911 4576 18368 4604
rect 17911 4573 17923 4576
rect 17865 4567 17923 4573
rect 18690 4564 18696 4616
rect 18748 4604 18754 4616
rect 18785 4607 18843 4613
rect 18785 4604 18797 4607
rect 18748 4576 18797 4604
rect 18748 4564 18754 4576
rect 18785 4573 18797 4576
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 19150 4564 19156 4616
rect 19208 4604 19214 4616
rect 19613 4607 19671 4613
rect 19613 4604 19625 4607
rect 19208 4576 19625 4604
rect 19208 4564 19214 4576
rect 19613 4573 19625 4576
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 20349 4607 20407 4613
rect 20349 4573 20361 4607
rect 20395 4604 20407 4607
rect 20958 4607 21016 4613
rect 20958 4604 20970 4607
rect 20395 4576 20970 4604
rect 20395 4573 20407 4576
rect 20349 4567 20407 4573
rect 20958 4573 20970 4576
rect 21004 4604 21016 4607
rect 21004 4576 21864 4604
rect 21004 4573 21016 4576
rect 20958 4567 21016 4573
rect 15160 4508 15608 4536
rect 15160 4496 15166 4508
rect 16942 4496 16948 4548
rect 17000 4496 17006 4548
rect 17129 4539 17187 4545
rect 17129 4505 17141 4539
rect 17175 4505 17187 4539
rect 17129 4499 17187 4505
rect 18509 4539 18567 4545
rect 18509 4505 18521 4539
rect 18555 4536 18567 4539
rect 18601 4539 18659 4545
rect 18601 4536 18613 4539
rect 18555 4508 18613 4536
rect 18555 4505 18567 4508
rect 18509 4499 18567 4505
rect 18601 4505 18613 4508
rect 18647 4505 18659 4539
rect 18601 4499 18659 4505
rect 14921 4471 14979 4477
rect 14921 4437 14933 4471
rect 14967 4437 14979 4471
rect 14921 4431 14979 4437
rect 15470 4428 15476 4480
rect 15528 4468 15534 4480
rect 15933 4471 15991 4477
rect 15933 4468 15945 4471
rect 15528 4440 15945 4468
rect 15528 4428 15534 4440
rect 15933 4437 15945 4440
rect 15979 4437 15991 4471
rect 15933 4431 15991 4437
rect 16485 4471 16543 4477
rect 16485 4437 16497 4471
rect 16531 4468 16543 4471
rect 17144 4468 17172 4499
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 19429 4539 19487 4545
rect 19429 4536 19441 4539
rect 19392 4508 19441 4536
rect 19392 4496 19398 4508
rect 19429 4505 19441 4508
rect 19475 4505 19487 4539
rect 19429 4499 19487 4505
rect 16531 4440 17172 4468
rect 19444 4468 19472 4499
rect 21836 4477 21864 4576
rect 22002 4564 22008 4616
rect 22060 4564 22066 4616
rect 19981 4471 20039 4477
rect 19981 4468 19993 4471
rect 19444 4440 19993 4468
rect 16531 4437 16543 4440
rect 16485 4431 16543 4437
rect 19981 4437 19993 4440
rect 20027 4437 20039 4471
rect 19981 4431 20039 4437
rect 20441 4471 20499 4477
rect 20441 4437 20453 4471
rect 20487 4468 20499 4471
rect 20855 4471 20913 4477
rect 20855 4468 20867 4471
rect 20487 4440 20867 4468
rect 20487 4437 20499 4440
rect 20441 4431 20499 4437
rect 20855 4437 20867 4440
rect 20901 4437 20913 4471
rect 20855 4431 20913 4437
rect 21821 4471 21879 4477
rect 21821 4437 21833 4471
rect 21867 4437 21879 4471
rect 21821 4431 21879 4437
rect 1104 4378 22356 4400
rect 1104 4326 4266 4378
rect 4318 4326 4330 4378
rect 4382 4326 4394 4378
rect 4446 4326 4458 4378
rect 4510 4326 4522 4378
rect 4574 4326 9579 4378
rect 9631 4326 9643 4378
rect 9695 4326 9707 4378
rect 9759 4326 9771 4378
rect 9823 4326 9835 4378
rect 9887 4326 14892 4378
rect 14944 4326 14956 4378
rect 15008 4326 15020 4378
rect 15072 4326 15084 4378
rect 15136 4326 15148 4378
rect 15200 4326 20205 4378
rect 20257 4326 20269 4378
rect 20321 4326 20333 4378
rect 20385 4326 20397 4378
rect 20449 4326 20461 4378
rect 20513 4326 22356 4378
rect 1104 4304 22356 4326
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 4065 4267 4123 4273
rect 4065 4264 4077 4267
rect 4028 4236 4077 4264
rect 4028 4224 4034 4236
rect 4065 4233 4077 4236
rect 4111 4233 4123 4267
rect 4065 4227 4123 4233
rect 7466 4224 7472 4276
rect 7524 4224 7530 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10045 4267 10103 4273
rect 10045 4264 10057 4267
rect 10008 4236 10057 4264
rect 10008 4224 10014 4236
rect 10045 4233 10057 4236
rect 10091 4233 10103 4267
rect 10045 4227 10103 4233
rect 10134 4224 10140 4276
rect 10192 4224 10198 4276
rect 13265 4267 13323 4273
rect 13265 4233 13277 4267
rect 13311 4264 13323 4267
rect 13538 4264 13544 4276
rect 13311 4236 13544 4264
rect 13311 4233 13323 4236
rect 13265 4227 13323 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 14369 4267 14427 4273
rect 14369 4264 14381 4267
rect 13872 4236 14381 4264
rect 13872 4224 13878 4236
rect 14369 4233 14381 4236
rect 14415 4233 14427 4267
rect 14369 4227 14427 4233
rect 18785 4267 18843 4273
rect 18785 4233 18797 4267
rect 18831 4264 18843 4267
rect 19058 4264 19064 4276
rect 18831 4236 19064 4264
rect 18831 4233 18843 4236
rect 18785 4227 18843 4233
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4196 4491 4199
rect 4798 4196 4804 4208
rect 4479 4168 4804 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 4798 4156 4804 4168
rect 4856 4196 4862 4208
rect 4856 4168 5120 4196
rect 4856 4156 4862 4168
rect 4890 4088 4896 4140
rect 4948 4088 4954 4140
rect 5092 4128 5120 4168
rect 5626 4156 5632 4208
rect 5684 4196 5690 4208
rect 5721 4199 5779 4205
rect 5721 4196 5733 4199
rect 5684 4168 5733 4196
rect 5684 4156 5690 4168
rect 5721 4165 5733 4168
rect 5767 4196 5779 4199
rect 6270 4196 6276 4208
rect 5767 4168 6276 4196
rect 5767 4165 5779 4168
rect 5721 4159 5779 4165
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 17218 4196 17224 4208
rect 15488 4168 17224 4196
rect 15488 4140 15516 4168
rect 17218 4156 17224 4168
rect 17276 4196 17282 4208
rect 19153 4199 19211 4205
rect 17276 4168 17356 4196
rect 17276 4156 17282 4168
rect 6114 4131 6172 4137
rect 6114 4128 6126 4131
rect 5092 4100 6126 4128
rect 6114 4097 6126 4100
rect 6160 4097 6172 4131
rect 6114 4091 6172 4097
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 7006 4128 7012 4140
rect 6696 4100 7012 4128
rect 6696 4088 6702 4100
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9456 4100 9689 4128
rect 9456 4088 9462 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 9907 4100 10364 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 4525 4063 4583 4069
rect 4525 4029 4537 4063
rect 4571 4029 4583 4063
rect 4525 4023 4583 4029
rect 4540 3992 4568 4023
rect 4706 4020 4712 4072
rect 4764 4020 4770 4072
rect 6733 4063 6791 4069
rect 6733 4029 6745 4063
rect 6779 4060 6791 4063
rect 6914 4060 6920 4072
rect 6779 4032 6920 4060
rect 6779 4029 6791 4032
rect 6733 4023 6791 4029
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7190 4020 7196 4072
rect 7248 4020 7254 4072
rect 7374 4020 7380 4072
rect 7432 4020 7438 4072
rect 6043 3995 6101 4001
rect 6043 3992 6055 3995
rect 4540 3964 6055 3992
rect 6043 3961 6055 3964
rect 6089 3961 6101 3995
rect 6043 3955 6101 3961
rect 7009 3995 7067 4001
rect 7009 3961 7021 3995
rect 7055 3992 7067 3995
rect 7282 3992 7288 4004
rect 7055 3964 7288 3992
rect 7055 3961 7067 3964
rect 7009 3955 7067 3961
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 7837 3995 7895 4001
rect 7837 3992 7849 3995
rect 7708 3964 7849 3992
rect 7708 3952 7714 3964
rect 7837 3961 7849 3964
rect 7883 3961 7895 3995
rect 9692 3992 9720 4091
rect 10336 4069 10364 4100
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 13538 4128 13544 4140
rect 12912 4100 13544 4128
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10367 4032 10824 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10796 4004 10824 4032
rect 11974 4020 11980 4072
rect 12032 4020 12038 4072
rect 12912 4069 12940 4100
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 13998 4088 14004 4140
rect 14056 4128 14062 4140
rect 15470 4128 15476 4140
rect 14056 4100 15476 4128
rect 14056 4088 14062 4100
rect 12069 4063 12127 4069
rect 12069 4029 12081 4063
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 13630 4060 13636 4072
rect 13127 4032 13636 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 10505 3995 10563 4001
rect 10505 3992 10517 3995
rect 9692 3964 10517 3992
rect 7837 3955 7895 3961
rect 10505 3961 10517 3964
rect 10551 3961 10563 3995
rect 10505 3955 10563 3961
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 10836 3964 11529 3992
rect 10836 3952 10842 3964
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 12084 3992 12112 4023
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 14108 4069 14136 4100
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 15657 4131 15715 4137
rect 15657 4097 15669 4131
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 16114 4128 16120 4140
rect 15887 4100 16120 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 14277 4063 14335 4069
rect 14277 4029 14289 4063
rect 14323 4029 14335 4063
rect 15672 4060 15700 4091
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 17034 4088 17040 4140
rect 17092 4088 17098 4140
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 15672 4032 16221 4060
rect 14277 4023 14335 4029
rect 16209 4029 16221 4032
rect 16255 4060 16267 4063
rect 16390 4060 16396 4072
rect 16255 4032 16396 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 11517 3955 11575 3961
rect 12059 3964 12112 3992
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 11054 3924 11060 3936
rect 7800 3896 11060 3924
rect 7800 3884 7806 3896
rect 11054 3884 11060 3896
rect 11112 3924 11118 3936
rect 12059 3924 12087 3964
rect 13998 3952 14004 4004
rect 14056 3992 14062 4004
rect 14292 3992 14320 4023
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16485 4063 16543 4069
rect 16485 4029 16497 4063
rect 16531 4060 16543 4063
rect 16666 4060 16672 4072
rect 16531 4032 16672 4060
rect 16531 4029 16543 4032
rect 16485 4023 16543 4029
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 17328 4069 17356 4168
rect 19153 4165 19165 4199
rect 19199 4196 19211 4199
rect 19426 4196 19432 4208
rect 19199 4168 19432 4196
rect 19199 4165 19211 4168
rect 19153 4159 19211 4165
rect 19426 4156 19432 4168
rect 19484 4156 19490 4208
rect 17129 4063 17187 4069
rect 17129 4029 17141 4063
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 14056 3964 14320 3992
rect 14056 3952 14062 3964
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 14737 3995 14795 4001
rect 14737 3992 14749 3995
rect 14608 3964 14749 3992
rect 14608 3952 14614 3964
rect 14737 3961 14749 3964
rect 14783 3961 14795 3995
rect 14737 3955 14795 3961
rect 15473 3995 15531 4001
rect 15473 3961 15485 3995
rect 15519 3992 15531 3995
rect 17144 3992 17172 4023
rect 19242 4020 19248 4072
rect 19300 4020 19306 4072
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19429 4063 19487 4069
rect 19429 4060 19441 4063
rect 19392 4032 19441 4060
rect 19392 4020 19398 4032
rect 19429 4029 19441 4032
rect 19475 4060 19487 4063
rect 19978 4060 19984 4072
rect 19475 4032 19984 4060
rect 19475 4029 19487 4032
rect 19429 4023 19487 4029
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 15519 3964 17172 3992
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 11112 3896 12087 3924
rect 13909 3927 13967 3933
rect 11112 3884 11118 3896
rect 13909 3893 13921 3927
rect 13955 3924 13967 3927
rect 14090 3924 14096 3936
rect 13955 3896 14096 3924
rect 13955 3893 13967 3896
rect 13909 3887 13967 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 16632 3896 16681 3924
rect 16632 3884 16638 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 1104 3834 22356 3856
rect 1104 3782 3606 3834
rect 3658 3782 3670 3834
rect 3722 3782 3734 3834
rect 3786 3782 3798 3834
rect 3850 3782 3862 3834
rect 3914 3782 8919 3834
rect 8971 3782 8983 3834
rect 9035 3782 9047 3834
rect 9099 3782 9111 3834
rect 9163 3782 9175 3834
rect 9227 3782 14232 3834
rect 14284 3782 14296 3834
rect 14348 3782 14360 3834
rect 14412 3782 14424 3834
rect 14476 3782 14488 3834
rect 14540 3782 19545 3834
rect 19597 3782 19609 3834
rect 19661 3782 19673 3834
rect 19725 3782 19737 3834
rect 19789 3782 19801 3834
rect 19853 3782 22356 3834
rect 1104 3760 22356 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 4890 3720 4896 3732
rect 1627 3692 4896 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5813 3723 5871 3729
rect 5813 3689 5825 3723
rect 5859 3720 5871 3723
rect 6822 3720 6828 3732
rect 5859 3692 6828 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7374 3680 7380 3732
rect 7432 3680 7438 3732
rect 9398 3680 9404 3732
rect 9456 3680 9462 3732
rect 11471 3723 11529 3729
rect 11471 3689 11483 3723
rect 11517 3720 11529 3723
rect 11974 3720 11980 3732
rect 11517 3692 11980 3720
rect 11517 3689 11529 3692
rect 11471 3683 11529 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 13449 3723 13507 3729
rect 13449 3689 13461 3723
rect 13495 3720 13507 3723
rect 13814 3720 13820 3732
rect 13495 3692 13820 3720
rect 13495 3689 13507 3692
rect 13449 3683 13507 3689
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 13998 3720 14004 3732
rect 13955 3692 14004 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 16577 3723 16635 3729
rect 16577 3689 16589 3723
rect 16623 3720 16635 3723
rect 16942 3720 16948 3732
rect 16623 3692 16948 3720
rect 16623 3689 16635 3692
rect 16577 3683 16635 3689
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 17034 3680 17040 3732
rect 17092 3680 17098 3732
rect 19242 3680 19248 3732
rect 19300 3729 19306 3732
rect 19300 3723 19349 3729
rect 19300 3689 19303 3723
rect 19337 3689 19349 3723
rect 19300 3683 19349 3689
rect 19300 3680 19306 3683
rect 6914 3652 6920 3664
rect 6012 3624 6920 3652
rect 6012 3593 6040 3624
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7024 3624 14780 3652
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 842 3408 848 3460
rect 900 3448 906 3460
rect 1489 3451 1547 3457
rect 1489 3448 1501 3451
rect 900 3420 1501 3448
rect 900 3408 906 3420
rect 1489 3417 1501 3420
rect 1535 3417 1547 3451
rect 6196 3448 6224 3547
rect 6270 3544 6276 3596
rect 6328 3584 6334 3596
rect 7024 3584 7052 3624
rect 6328 3556 7052 3584
rect 6328 3544 6334 3556
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 7558 3584 7564 3596
rect 7340 3556 7564 3584
rect 7340 3544 7346 3556
rect 7558 3544 7564 3556
rect 7616 3584 7622 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 7616 3556 10057 3584
rect 7616 3544 7622 3556
rect 10045 3553 10057 3556
rect 10091 3584 10103 3587
rect 10594 3584 10600 3596
rect 10091 3556 10600 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 13081 3587 13139 3593
rect 13081 3553 13093 3587
rect 13127 3553 13139 3587
rect 13081 3547 13139 3553
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7193 3519 7251 3525
rect 7193 3516 7205 3519
rect 6972 3488 7205 3516
rect 6972 3476 6978 3488
rect 7193 3485 7205 3488
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 11400 3519 11458 3525
rect 11400 3516 11412 3519
rect 11296 3488 11412 3516
rect 11296 3476 11302 3488
rect 11400 3485 11412 3488
rect 11446 3516 11458 3519
rect 11882 3516 11888 3528
rect 11446 3488 11888 3516
rect 11446 3485 11458 3488
rect 11400 3479 11458 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 6638 3448 6644 3460
rect 6196 3420 6644 3448
rect 1489 3411 1547 3417
rect 6638 3408 6644 3420
rect 6696 3448 6702 3460
rect 7009 3451 7067 3457
rect 7009 3448 7021 3451
rect 6696 3420 7021 3448
rect 6696 3408 6702 3420
rect 7009 3417 7021 3420
rect 7055 3417 7067 3451
rect 7009 3411 7067 3417
rect 9769 3451 9827 3457
rect 9769 3417 9781 3451
rect 9815 3448 9827 3451
rect 10042 3448 10048 3460
rect 9815 3420 10048 3448
rect 9815 3417 9827 3420
rect 9769 3411 9827 3417
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 13096 3448 13124 3547
rect 13265 3519 13323 3525
rect 13265 3485 13277 3519
rect 13311 3516 13323 3519
rect 13630 3516 13636 3528
rect 13311 3488 13636 3516
rect 13311 3485 13323 3488
rect 13265 3479 13323 3485
rect 13630 3476 13636 3488
rect 13688 3516 13694 3528
rect 13688 3488 13768 3516
rect 13688 3476 13694 3488
rect 13538 3448 13544 3460
rect 13096 3420 13544 3448
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 13740 3457 13768 3488
rect 14182 3476 14188 3528
rect 14240 3525 14246 3528
rect 14240 3519 14268 3525
rect 14256 3485 14268 3519
rect 14240 3479 14268 3485
rect 14240 3476 14246 3479
rect 13725 3451 13783 3457
rect 13725 3417 13737 3451
rect 13771 3448 13783 3451
rect 14642 3448 14648 3460
rect 13771 3420 14648 3448
rect 13771 3417 13783 3420
rect 13725 3411 13783 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 14752 3457 14780 3624
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16209 3587 16267 3593
rect 16209 3584 16221 3587
rect 16172 3556 16221 3584
rect 16172 3544 16178 3556
rect 16209 3553 16221 3556
rect 16255 3584 16267 3587
rect 16482 3584 16488 3596
rect 16255 3556 16488 3584
rect 16255 3553 16267 3556
rect 16209 3547 16267 3553
rect 16482 3544 16488 3556
rect 16540 3584 16546 3596
rect 16669 3587 16727 3593
rect 16669 3584 16681 3587
rect 16540 3556 16681 3584
rect 16540 3544 16546 3556
rect 16669 3553 16681 3556
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 16390 3476 16396 3528
rect 16448 3516 16454 3528
rect 16850 3516 16856 3528
rect 16448 3488 16856 3516
rect 16448 3476 16454 3488
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 17196 3519 17254 3525
rect 17196 3485 17208 3519
rect 17242 3516 17254 3519
rect 17310 3516 17316 3528
rect 17242 3488 17316 3516
rect 17242 3485 17254 3488
rect 17196 3479 17254 3485
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 19426 3525 19432 3528
rect 19394 3519 19432 3525
rect 19394 3485 19406 3519
rect 19394 3479 19432 3485
rect 19426 3476 19432 3479
rect 19484 3476 19490 3528
rect 14737 3451 14795 3457
rect 14737 3417 14749 3451
rect 14783 3448 14795 3451
rect 17034 3448 17040 3460
rect 14783 3420 17040 3448
rect 14783 3417 14795 3420
rect 14737 3411 14795 3417
rect 17034 3408 17040 3420
rect 17092 3408 17098 3460
rect 9861 3383 9919 3389
rect 9861 3349 9873 3383
rect 9907 3380 9919 3383
rect 9950 3380 9956 3392
rect 9907 3352 9956 3380
rect 9907 3349 9919 3352
rect 9861 3343 9919 3349
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 14139 3383 14197 3389
rect 14139 3349 14151 3383
rect 14185 3380 14197 3383
rect 14274 3380 14280 3392
rect 14185 3352 14280 3380
rect 14185 3349 14197 3352
rect 14139 3343 14197 3349
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 14461 3383 14519 3389
rect 14461 3349 14473 3383
rect 14507 3380 14519 3383
rect 15286 3380 15292 3392
rect 14507 3352 15292 3380
rect 14507 3349 14519 3352
rect 14461 3343 14519 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 17267 3383 17325 3389
rect 17267 3349 17279 3383
rect 17313 3380 17325 3383
rect 17862 3380 17868 3392
rect 17313 3352 17868 3380
rect 17313 3349 17325 3352
rect 17267 3343 17325 3349
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 1104 3290 22356 3312
rect 1104 3238 4266 3290
rect 4318 3238 4330 3290
rect 4382 3238 4394 3290
rect 4446 3238 4458 3290
rect 4510 3238 4522 3290
rect 4574 3238 9579 3290
rect 9631 3238 9643 3290
rect 9695 3238 9707 3290
rect 9759 3238 9771 3290
rect 9823 3238 9835 3290
rect 9887 3238 14892 3290
rect 14944 3238 14956 3290
rect 15008 3238 15020 3290
rect 15072 3238 15084 3290
rect 15136 3238 15148 3290
rect 15200 3238 20205 3290
rect 20257 3238 20269 3290
rect 20321 3238 20333 3290
rect 20385 3238 20397 3290
rect 20449 3238 20461 3290
rect 20513 3238 22356 3290
rect 1104 3216 22356 3238
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6972 3148 7113 3176
rect 6972 3136 6978 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 9815 3179 9873 3185
rect 9815 3145 9827 3179
rect 9861 3176 9873 3179
rect 9950 3176 9956 3188
rect 9861 3148 9956 3176
rect 9861 3145 9873 3148
rect 9815 3139 9873 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13596 3148 13829 3176
rect 13596 3136 13602 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 13817 3139 13875 3145
rect 14274 3136 14280 3188
rect 14332 3136 14338 3188
rect 14642 3136 14648 3188
rect 14700 3136 14706 3188
rect 16482 3136 16488 3188
rect 16540 3176 16546 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 16540 3148 16681 3176
rect 16540 3136 16546 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 16669 3139 16727 3145
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 16908 3148 17509 3176
rect 16908 3136 16914 3148
rect 17497 3145 17509 3148
rect 17543 3145 17555 3179
rect 17497 3139 17555 3145
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 17957 3179 18015 3185
rect 17957 3176 17969 3179
rect 17920 3148 17969 3176
rect 17920 3136 17926 3148
rect 17957 3145 17969 3148
rect 18003 3145 18015 3179
rect 17957 3139 18015 3145
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 5592 3080 7481 3108
rect 5592 3068 5598 3080
rect 7469 3077 7481 3080
rect 7515 3108 7527 3111
rect 19334 3108 19340 3120
rect 7515 3080 8156 3108
rect 7515 3077 7527 3080
rect 7469 3071 7527 3077
rect 6914 3049 6920 3052
rect 6892 3043 6920 3049
rect 6892 3009 6904 3043
rect 6892 3003 6920 3009
rect 6914 3000 6920 3003
rect 6972 3000 6978 3052
rect 8128 3049 8156 3080
rect 14476 3080 19340 3108
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7975 3043 8033 3049
rect 7975 3040 7987 3043
rect 7607 3012 7987 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7975 3009 7987 3012
rect 8021 3009 8033 3043
rect 7975 3003 8033 3009
rect 8078 3043 8156 3049
rect 8078 3009 8090 3043
rect 8124 3012 8156 3043
rect 9918 3043 9976 3049
rect 8124 3009 8136 3012
rect 8078 3003 8136 3009
rect 9918 3009 9930 3043
rect 9964 3040 9976 3043
rect 10042 3040 10048 3052
rect 9964 3012 10048 3040
rect 9964 3009 9976 3012
rect 9918 3003 9976 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 13608 3043 13666 3049
rect 13608 3009 13620 3043
rect 13654 3040 13666 3043
rect 13814 3040 13820 3052
rect 13654 3012 13820 3040
rect 13654 3009 13666 3012
rect 13608 3003 13666 3009
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 14182 3000 14188 3052
rect 14240 3000 14246 3052
rect 7742 2932 7748 2984
rect 7800 2932 7806 2984
rect 14476 2981 14504 3080
rect 15010 3000 15016 3052
rect 15068 3000 15074 3052
rect 16352 3043 16410 3049
rect 16352 3009 16364 3043
rect 16398 3040 16410 3043
rect 17034 3040 17040 3052
rect 16398 3012 17040 3040
rect 16398 3009 16410 3012
rect 16352 3003 16410 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 15105 2975 15163 2981
rect 15105 2941 15117 2975
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 13679 2907 13737 2913
rect 13679 2873 13691 2907
rect 13725 2904 13737 2907
rect 15120 2904 15148 2935
rect 15286 2932 15292 2984
rect 15344 2932 15350 2984
rect 17236 2981 17264 3080
rect 19334 3068 19340 3080
rect 19392 3068 19398 3120
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 17865 3043 17923 3049
rect 17865 3040 17877 3043
rect 17368 3012 17877 3040
rect 17368 3000 17374 3012
rect 17865 3009 17877 3012
rect 17911 3040 17923 3043
rect 20070 3040 20076 3052
rect 17911 3012 20076 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 16439 2975 16497 2981
rect 16439 2941 16451 2975
rect 16485 2972 16497 2975
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 16485 2944 17141 2972
rect 16485 2941 16497 2944
rect 16439 2935 16497 2941
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2972 18199 2975
rect 20622 2972 20628 2984
rect 18187 2944 20628 2972
rect 18187 2941 18199 2944
rect 18141 2935 18199 2941
rect 13725 2876 15148 2904
rect 15304 2904 15332 2932
rect 18156 2904 18184 2935
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 15304 2876 18184 2904
rect 13725 2873 13737 2876
rect 13679 2867 13737 2873
rect 7006 2845 7012 2848
rect 6963 2839 7012 2845
rect 6963 2805 6975 2839
rect 7009 2805 7012 2839
rect 6963 2799 7012 2805
rect 7006 2796 7012 2799
rect 7064 2796 7070 2848
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 14918 2836 14924 2848
rect 14240 2808 14924 2836
rect 14240 2796 14246 2808
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 1104 2746 22356 2768
rect 1104 2694 3606 2746
rect 3658 2694 3670 2746
rect 3722 2694 3734 2746
rect 3786 2694 3798 2746
rect 3850 2694 3862 2746
rect 3914 2694 8919 2746
rect 8971 2694 8983 2746
rect 9035 2694 9047 2746
rect 9099 2694 9111 2746
rect 9163 2694 9175 2746
rect 9227 2694 14232 2746
rect 14284 2694 14296 2746
rect 14348 2694 14360 2746
rect 14412 2694 14424 2746
rect 14476 2694 14488 2746
rect 14540 2694 19545 2746
rect 19597 2694 19609 2746
rect 19661 2694 19673 2746
rect 19725 2694 19737 2746
rect 19789 2694 19801 2746
rect 19853 2694 22356 2746
rect 1104 2672 22356 2694
rect 4798 2592 4804 2644
rect 4856 2592 4862 2644
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 5534 2632 5540 2644
rect 5491 2604 5540 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 6914 2632 6920 2644
rect 6595 2604 6920 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10042 2632 10048 2644
rect 9999 2604 10048 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10410 2592 10416 2644
rect 10468 2592 10474 2644
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11572 2604 11713 2632
rect 11572 2592 11578 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 12526 2592 12532 2644
rect 12584 2592 12590 2644
rect 14918 2592 14924 2644
rect 14976 2592 14982 2644
rect 17034 2592 17040 2644
rect 17092 2632 17098 2644
rect 18141 2635 18199 2641
rect 18141 2632 18153 2635
rect 17092 2604 18153 2632
rect 17092 2592 17098 2604
rect 18141 2601 18153 2604
rect 18187 2601 18199 2635
rect 18141 2595 18199 2601
rect 19426 2592 19432 2644
rect 19484 2592 19490 2644
rect 20070 2592 20076 2644
rect 20128 2592 20134 2644
rect 3513 2567 3571 2573
rect 3513 2533 3525 2567
rect 3559 2533 3571 2567
rect 3513 2527 3571 2533
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 9309 2567 9367 2573
rect 4203 2536 9260 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 3528 2496 3556 2527
rect 3528 2468 6914 2496
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3292 2400 3341 2428
rect 3292 2388 3298 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 5224 2400 5273 2428
rect 5224 2388 5230 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 6454 2428 6460 2440
rect 6411 2400 6460 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 6196 2360 6224 2391
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 6886 2428 6914 2468
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 7064 2468 7113 2496
rect 7064 2456 7070 2468
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 7101 2459 7159 2465
rect 7282 2456 7288 2508
rect 7340 2456 7346 2508
rect 6886 2400 7420 2428
rect 6196 2332 6776 2360
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 5997 2295 6055 2301
rect 5997 2292 6009 2295
rect 5868 2264 6009 2292
rect 5868 2252 5874 2264
rect 5997 2261 6009 2264
rect 6043 2261 6055 2295
rect 5997 2255 6055 2261
rect 6638 2252 6644 2304
rect 6696 2252 6702 2304
rect 6748 2292 6776 2332
rect 6914 2320 6920 2372
rect 6972 2360 6978 2372
rect 7009 2363 7067 2369
rect 7009 2360 7021 2363
rect 6972 2332 7021 2360
rect 6972 2320 6978 2332
rect 7009 2329 7021 2332
rect 7055 2329 7067 2363
rect 7282 2360 7288 2372
rect 7009 2323 7067 2329
rect 7116 2332 7288 2360
rect 7116 2292 7144 2332
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 7392 2360 7420 2400
rect 7466 2388 7472 2440
rect 7524 2388 7530 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8570 2428 8576 2440
rect 8527 2400 8576 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9232 2360 9260 2536
rect 9309 2533 9321 2567
rect 9355 2564 9367 2567
rect 11330 2564 11336 2576
rect 9355 2536 11336 2564
rect 9355 2533 9367 2536
rect 9309 2527 9367 2533
rect 11330 2524 11336 2536
rect 11388 2524 11394 2576
rect 12066 2524 12072 2576
rect 12124 2564 12130 2576
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 12124 2536 13645 2564
rect 12124 2524 12130 2536
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 13633 2527 13691 2533
rect 13814 2524 13820 2576
rect 13872 2564 13878 2576
rect 15010 2564 15016 2576
rect 13872 2536 15016 2564
rect 13872 2524 13878 2536
rect 15010 2524 15016 2536
rect 15068 2564 15074 2576
rect 17497 2567 17555 2573
rect 17497 2564 17509 2567
rect 15068 2536 17509 2564
rect 15068 2524 15074 2536
rect 17497 2533 17509 2536
rect 17543 2533 17555 2567
rect 17497 2527 17555 2533
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 9950 2428 9956 2440
rect 9815 2400 9956 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 11020 2400 11069 2428
rect 11020 2388 11026 2400
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11664 2400 11897 2428
rect 11664 2388 11670 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2428 13047 2431
rect 13078 2428 13084 2440
rect 13035 2400 13084 2428
rect 13035 2397 13047 2400
rect 12989 2391 13047 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 13817 2431 13875 2437
rect 13817 2428 13829 2431
rect 13596 2400 13829 2428
rect 13596 2388 13602 2400
rect 13817 2397 13829 2400
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13964 2400 14289 2428
rect 13964 2388 13970 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 14792 2400 15117 2428
rect 14792 2388 14798 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15562 2388 15568 2440
rect 15620 2388 15626 2440
rect 16206 2388 16212 2440
rect 16264 2388 16270 2440
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17460 2400 17693 2428
rect 17460 2388 17466 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18104 2400 18337 2428
rect 18104 2388 18110 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 20036 2400 20269 2428
rect 20036 2388 20042 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 11790 2360 11796 2372
rect 7392 2332 8800 2360
rect 9232 2332 11796 2360
rect 6748 2264 7144 2292
rect 7190 2252 7196 2304
rect 7248 2292 7254 2304
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 7248 2264 7665 2292
rect 7248 2252 7254 2264
rect 7653 2261 7665 2264
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8444 2264 8677 2292
rect 8444 2252 8450 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8772 2292 8800 2332
rect 11790 2320 11796 2332
rect 11848 2320 11854 2372
rect 12894 2320 12900 2372
rect 12952 2360 12958 2372
rect 13265 2363 13323 2369
rect 13265 2360 13277 2363
rect 12952 2332 13277 2360
rect 12952 2320 12958 2332
rect 13265 2329 13277 2332
rect 13311 2329 13323 2363
rect 13265 2323 13323 2329
rect 11146 2292 11152 2304
rect 8772 2264 11152 2292
rect 8665 2255 8723 2261
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 14240 2264 14473 2292
rect 14240 2252 14246 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15528 2264 15761 2292
rect 15528 2252 15534 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16393 2295 16451 2301
rect 16393 2292 16405 2295
rect 16172 2264 16405 2292
rect 16172 2252 16178 2264
rect 16393 2261 16405 2264
rect 16439 2261 16451 2295
rect 16393 2255 16451 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18969 2295 19027 2301
rect 18969 2292 18981 2295
rect 18748 2264 18981 2292
rect 18748 2252 18754 2264
rect 18969 2261 18981 2264
rect 19015 2261 19027 2295
rect 18969 2255 19027 2261
rect 1104 2202 22356 2224
rect 1104 2150 4266 2202
rect 4318 2150 4330 2202
rect 4382 2150 4394 2202
rect 4446 2150 4458 2202
rect 4510 2150 4522 2202
rect 4574 2150 9579 2202
rect 9631 2150 9643 2202
rect 9695 2150 9707 2202
rect 9759 2150 9771 2202
rect 9823 2150 9835 2202
rect 9887 2150 14892 2202
rect 14944 2150 14956 2202
rect 15008 2150 15020 2202
rect 15072 2150 15084 2202
rect 15136 2150 15148 2202
rect 15200 2150 20205 2202
rect 20257 2150 20269 2202
rect 20321 2150 20333 2202
rect 20385 2150 20397 2202
rect 20449 2150 20461 2202
rect 20513 2150 22356 2202
rect 1104 2128 22356 2150
<< via1 >>
rect 3606 23366 3658 23418
rect 3670 23366 3722 23418
rect 3734 23366 3786 23418
rect 3798 23366 3850 23418
rect 3862 23366 3914 23418
rect 8919 23366 8971 23418
rect 8983 23366 9035 23418
rect 9047 23366 9099 23418
rect 9111 23366 9163 23418
rect 9175 23366 9227 23418
rect 14232 23366 14284 23418
rect 14296 23366 14348 23418
rect 14360 23366 14412 23418
rect 14424 23366 14476 23418
rect 14488 23366 14540 23418
rect 19545 23366 19597 23418
rect 19609 23366 19661 23418
rect 19673 23366 19725 23418
rect 19737 23366 19789 23418
rect 19801 23366 19853 23418
rect 7104 23264 7156 23316
rect 8024 23307 8076 23316
rect 8024 23273 8033 23307
rect 8033 23273 8067 23307
rect 8067 23273 8076 23307
rect 8024 23264 8076 23273
rect 11612 23307 11664 23316
rect 11612 23273 11621 23307
rect 11621 23273 11655 23307
rect 11655 23273 11664 23307
rect 11612 23264 11664 23273
rect 14096 23264 14148 23316
rect 16764 23264 16816 23316
rect 18328 23307 18380 23316
rect 18328 23273 18337 23307
rect 18337 23273 18371 23307
rect 18371 23273 18380 23307
rect 18328 23264 18380 23273
rect 11060 23196 11112 23248
rect 12256 23239 12308 23248
rect 12256 23205 12265 23239
rect 12265 23205 12299 23239
rect 12299 23205 12308 23239
rect 12256 23196 12308 23205
rect 16120 23196 16172 23248
rect 4804 23103 4856 23112
rect 4804 23069 4813 23103
rect 4813 23069 4847 23103
rect 4847 23069 4856 23103
rect 4804 23060 4856 23069
rect 5264 23103 5316 23112
rect 5264 23069 5273 23103
rect 5273 23069 5307 23103
rect 5307 23069 5316 23103
rect 5264 23060 5316 23069
rect 6552 23103 6604 23112
rect 6552 23069 6561 23103
rect 6561 23069 6595 23103
rect 6595 23069 6604 23103
rect 6552 23060 6604 23069
rect 8392 23060 8444 23112
rect 9312 23060 9364 23112
rect 9680 23060 9732 23112
rect 10416 23103 10468 23112
rect 10416 23069 10425 23103
rect 10425 23069 10459 23103
rect 10459 23069 10468 23103
rect 10416 23060 10468 23069
rect 10968 23060 11020 23112
rect 7288 23035 7340 23044
rect 7288 23001 7297 23035
rect 7297 23001 7331 23035
rect 7331 23001 7340 23035
rect 7288 22992 7340 23001
rect 7932 23035 7984 23044
rect 7932 23001 7941 23035
rect 7941 23001 7975 23035
rect 7975 23001 7984 23035
rect 7932 22992 7984 23001
rect 13360 23128 13412 23180
rect 12900 23060 12952 23112
rect 13544 23060 13596 23112
rect 15108 23103 15160 23112
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 15568 23103 15620 23112
rect 15568 23069 15577 23103
rect 15577 23069 15611 23103
rect 15611 23069 15620 23103
rect 15568 23060 15620 23069
rect 15660 23060 15712 23112
rect 17408 23060 17460 23112
rect 18972 23103 19024 23112
rect 18972 23069 18981 23103
rect 18981 23069 19015 23103
rect 19015 23069 19024 23103
rect 18972 23060 19024 23069
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 11888 23035 11940 23044
rect 11888 23001 11897 23035
rect 11897 23001 11931 23035
rect 11931 23001 11940 23035
rect 11888 22992 11940 23001
rect 12808 22992 12860 23044
rect 14004 22992 14056 23044
rect 16764 23035 16816 23044
rect 16764 23001 16773 23035
rect 16773 23001 16807 23035
rect 16807 23001 16816 23035
rect 16764 22992 16816 23001
rect 17316 23035 17368 23044
rect 17316 23001 17325 23035
rect 17325 23001 17359 23035
rect 17359 23001 17368 23035
rect 17316 22992 17368 23001
rect 18052 22992 18104 23044
rect 4620 22967 4672 22976
rect 4620 22933 4629 22967
rect 4629 22933 4663 22967
rect 4663 22933 4672 22967
rect 4620 22924 4672 22933
rect 5448 22967 5500 22976
rect 5448 22933 5457 22967
rect 5457 22933 5491 22967
rect 5491 22933 5500 22967
rect 5448 22924 5500 22933
rect 7748 22924 7800 22976
rect 8392 22924 8444 22976
rect 9956 22967 10008 22976
rect 9956 22933 9965 22967
rect 9965 22933 9999 22967
rect 9999 22933 10008 22967
rect 9956 22924 10008 22933
rect 10876 22924 10928 22976
rect 10968 22924 11020 22976
rect 11704 22924 11756 22976
rect 12624 22967 12676 22976
rect 12624 22933 12633 22967
rect 12633 22933 12667 22967
rect 12667 22933 12676 22967
rect 12624 22924 12676 22933
rect 13084 22967 13136 22976
rect 13084 22933 13093 22967
rect 13093 22933 13127 22967
rect 13127 22933 13136 22967
rect 13084 22924 13136 22933
rect 13636 22967 13688 22976
rect 13636 22933 13645 22967
rect 13645 22933 13679 22967
rect 13679 22933 13688 22967
rect 13636 22924 13688 22933
rect 13912 22967 13964 22976
rect 13912 22933 13921 22967
rect 13921 22933 13955 22967
rect 13955 22933 13964 22967
rect 13912 22924 13964 22933
rect 14556 22924 14608 22976
rect 15384 22967 15436 22976
rect 15384 22933 15393 22967
rect 15393 22933 15427 22967
rect 15427 22933 15436 22967
rect 15384 22924 15436 22933
rect 15752 22924 15804 22976
rect 16120 22967 16172 22976
rect 16120 22933 16129 22967
rect 16129 22933 16163 22967
rect 16163 22933 16172 22967
rect 16120 22924 16172 22933
rect 16488 22924 16540 22976
rect 19432 22924 19484 22976
rect 4266 22822 4318 22874
rect 4330 22822 4382 22874
rect 4394 22822 4446 22874
rect 4458 22822 4510 22874
rect 4522 22822 4574 22874
rect 9579 22822 9631 22874
rect 9643 22822 9695 22874
rect 9707 22822 9759 22874
rect 9771 22822 9823 22874
rect 9835 22822 9887 22874
rect 14892 22822 14944 22874
rect 14956 22822 15008 22874
rect 15020 22822 15072 22874
rect 15084 22822 15136 22874
rect 15148 22822 15200 22874
rect 20205 22822 20257 22874
rect 20269 22822 20321 22874
rect 20333 22822 20385 22874
rect 20397 22822 20449 22874
rect 20461 22822 20513 22874
rect 7748 22763 7800 22772
rect 7748 22729 7757 22763
rect 7757 22729 7791 22763
rect 7791 22729 7800 22763
rect 7748 22720 7800 22729
rect 848 22584 900 22636
rect 8392 22627 8444 22636
rect 8392 22593 8400 22627
rect 8400 22593 8444 22627
rect 8392 22584 8444 22593
rect 13084 22720 13136 22772
rect 16120 22720 16172 22772
rect 14096 22652 14148 22704
rect 2688 22516 2740 22568
rect 7012 22516 7064 22568
rect 10968 22516 11020 22568
rect 13360 22559 13412 22568
rect 13360 22525 13369 22559
rect 13369 22525 13403 22559
rect 13403 22525 13412 22559
rect 13360 22516 13412 22525
rect 13636 22627 13688 22636
rect 13636 22593 13670 22627
rect 13670 22593 13688 22627
rect 13636 22584 13688 22593
rect 15660 22584 15712 22636
rect 16488 22627 16540 22636
rect 16488 22593 16496 22627
rect 16496 22593 16540 22627
rect 16488 22584 16540 22593
rect 16672 22627 16724 22636
rect 16672 22593 16681 22627
rect 16681 22593 16715 22627
rect 16715 22593 16724 22627
rect 16672 22584 16724 22593
rect 13912 22516 13964 22568
rect 4896 22448 4948 22500
rect 7104 22380 7156 22432
rect 8300 22380 8352 22432
rect 12440 22380 12492 22432
rect 15476 22423 15528 22432
rect 15476 22389 15485 22423
rect 15485 22389 15519 22423
rect 15519 22389 15528 22423
rect 15476 22380 15528 22389
rect 16672 22380 16724 22432
rect 19892 22380 19944 22432
rect 3606 22278 3658 22330
rect 3670 22278 3722 22330
rect 3734 22278 3786 22330
rect 3798 22278 3850 22330
rect 3862 22278 3914 22330
rect 8919 22278 8971 22330
rect 8983 22278 9035 22330
rect 9047 22278 9099 22330
rect 9111 22278 9163 22330
rect 9175 22278 9227 22330
rect 14232 22278 14284 22330
rect 14296 22278 14348 22330
rect 14360 22278 14412 22330
rect 14424 22278 14476 22330
rect 14488 22278 14540 22330
rect 19545 22278 19597 22330
rect 19609 22278 19661 22330
rect 19673 22278 19725 22330
rect 19737 22278 19789 22330
rect 19801 22278 19853 22330
rect 848 21972 900 22024
rect 7104 22108 7156 22160
rect 7748 22040 7800 22092
rect 12624 22108 12676 22160
rect 8576 22083 8628 22092
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 8576 22040 8628 22049
rect 13268 22083 13320 22092
rect 13268 22049 13277 22083
rect 13277 22049 13311 22083
rect 13311 22049 13320 22083
rect 13268 22040 13320 22049
rect 13912 22040 13964 22092
rect 14096 22040 14148 22092
rect 15752 22108 15804 22160
rect 15476 22040 15528 22092
rect 15568 22083 15620 22092
rect 15568 22049 15577 22083
rect 15577 22049 15611 22083
rect 15611 22049 15620 22083
rect 15568 22040 15620 22049
rect 15660 22040 15712 22092
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 7380 21879 7432 21888
rect 7380 21845 7389 21879
rect 7389 21845 7423 21879
rect 7423 21845 7432 21879
rect 7380 21836 7432 21845
rect 8484 21972 8536 22024
rect 13728 22015 13780 22024
rect 13728 21981 13737 22015
rect 13737 21981 13771 22015
rect 13771 21981 13780 22015
rect 13728 21972 13780 21981
rect 12440 21947 12492 21956
rect 12440 21913 12449 21947
rect 12449 21913 12483 21947
rect 12483 21913 12492 21947
rect 12440 21904 12492 21913
rect 12624 21947 12676 21956
rect 12624 21913 12633 21947
rect 12633 21913 12667 21947
rect 12667 21913 12676 21947
rect 12624 21904 12676 21913
rect 12716 21879 12768 21888
rect 12716 21845 12725 21879
rect 12725 21845 12759 21879
rect 12759 21845 12768 21879
rect 12716 21836 12768 21845
rect 14648 21836 14700 21888
rect 15936 21836 15988 21888
rect 4266 21734 4318 21786
rect 4330 21734 4382 21786
rect 4394 21734 4446 21786
rect 4458 21734 4510 21786
rect 4522 21734 4574 21786
rect 9579 21734 9631 21786
rect 9643 21734 9695 21786
rect 9707 21734 9759 21786
rect 9771 21734 9823 21786
rect 9835 21734 9887 21786
rect 14892 21734 14944 21786
rect 14956 21734 15008 21786
rect 15020 21734 15072 21786
rect 15084 21734 15136 21786
rect 15148 21734 15200 21786
rect 20205 21734 20257 21786
rect 20269 21734 20321 21786
rect 20333 21734 20385 21786
rect 20397 21734 20449 21786
rect 20461 21734 20513 21786
rect 5448 21632 5500 21684
rect 8300 21632 8352 21684
rect 15936 21675 15988 21684
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 848 21496 900 21548
rect 4620 21496 4672 21548
rect 4160 21428 4212 21480
rect 7104 21539 7156 21548
rect 7104 21505 7113 21539
rect 7113 21505 7147 21539
rect 7147 21505 7156 21539
rect 7104 21496 7156 21505
rect 8024 21496 8076 21548
rect 4988 21360 5040 21412
rect 4528 21292 4580 21344
rect 5540 21292 5592 21344
rect 7196 21292 7248 21344
rect 15476 21564 15528 21616
rect 8484 21496 8536 21548
rect 12624 21496 12676 21548
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 12440 21428 12492 21480
rect 13728 21428 13780 21480
rect 15476 21471 15528 21480
rect 15476 21437 15485 21471
rect 15485 21437 15519 21471
rect 15519 21437 15528 21471
rect 15476 21428 15528 21437
rect 8576 21360 8628 21412
rect 12624 21360 12676 21412
rect 8300 21292 8352 21344
rect 13176 21335 13228 21344
rect 13176 21301 13185 21335
rect 13185 21301 13219 21335
rect 13219 21301 13228 21335
rect 13176 21292 13228 21301
rect 13452 21292 13504 21344
rect 15844 21335 15896 21344
rect 15844 21301 15853 21335
rect 15853 21301 15887 21335
rect 15887 21301 15896 21335
rect 15844 21292 15896 21301
rect 3606 21190 3658 21242
rect 3670 21190 3722 21242
rect 3734 21190 3786 21242
rect 3798 21190 3850 21242
rect 3862 21190 3914 21242
rect 8919 21190 8971 21242
rect 8983 21190 9035 21242
rect 9047 21190 9099 21242
rect 9111 21190 9163 21242
rect 9175 21190 9227 21242
rect 14232 21190 14284 21242
rect 14296 21190 14348 21242
rect 14360 21190 14412 21242
rect 14424 21190 14476 21242
rect 14488 21190 14540 21242
rect 19545 21190 19597 21242
rect 19609 21190 19661 21242
rect 19673 21190 19725 21242
rect 19737 21190 19789 21242
rect 19801 21190 19853 21242
rect 2688 21020 2740 21072
rect 4896 21020 4948 21072
rect 15660 21020 15712 21072
rect 4528 20995 4580 21004
rect 4528 20961 4537 20995
rect 4537 20961 4571 20995
rect 4571 20961 4580 20995
rect 4528 20952 4580 20961
rect 4712 20995 4764 21004
rect 4712 20961 4721 20995
rect 4721 20961 4755 20995
rect 4755 20961 4764 20995
rect 4712 20952 4764 20961
rect 6828 20952 6880 21004
rect 7196 20952 7248 21004
rect 4896 20927 4948 20936
rect 4896 20893 4905 20927
rect 4905 20893 4939 20927
rect 4939 20893 4948 20927
rect 4896 20884 4948 20893
rect 4620 20816 4672 20868
rect 4712 20816 4764 20868
rect 7012 20884 7064 20936
rect 7472 20927 7524 20936
rect 7472 20893 7481 20927
rect 7481 20893 7515 20927
rect 7515 20893 7524 20927
rect 7472 20884 7524 20893
rect 8300 20927 8352 20936
rect 8300 20893 8309 20927
rect 8309 20893 8343 20927
rect 8343 20893 8352 20927
rect 8300 20884 8352 20893
rect 13452 20927 13504 20936
rect 13452 20893 13461 20927
rect 13461 20893 13495 20927
rect 13495 20893 13504 20927
rect 13452 20884 13504 20893
rect 15292 20884 15344 20936
rect 17132 20884 17184 20936
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 18328 20884 18380 20936
rect 19892 20995 19944 21004
rect 19892 20961 19901 20995
rect 19901 20961 19935 20995
rect 19935 20961 19944 20995
rect 19892 20952 19944 20961
rect 20536 20952 20588 21004
rect 19432 20884 19484 20936
rect 22008 20927 22060 20936
rect 22008 20893 22017 20927
rect 22017 20893 22051 20927
rect 22051 20893 22060 20927
rect 22008 20884 22060 20893
rect 5540 20816 5592 20868
rect 5724 20816 5776 20868
rect 13636 20859 13688 20868
rect 13636 20825 13645 20859
rect 13645 20825 13679 20859
rect 13679 20825 13688 20859
rect 13636 20816 13688 20825
rect 15844 20816 15896 20868
rect 18604 20816 18656 20868
rect 19064 20859 19116 20868
rect 19064 20825 19073 20859
rect 19073 20825 19107 20859
rect 19107 20825 19116 20859
rect 19064 20816 19116 20825
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 3976 20748 4028 20800
rect 5448 20791 5500 20800
rect 5448 20757 5457 20791
rect 5457 20757 5491 20791
rect 5491 20757 5500 20791
rect 5448 20748 5500 20757
rect 9312 20748 9364 20800
rect 18236 20791 18288 20800
rect 18236 20757 18245 20791
rect 18245 20757 18279 20791
rect 18279 20757 18288 20791
rect 18236 20748 18288 20757
rect 18696 20791 18748 20800
rect 18696 20757 18705 20791
rect 18705 20757 18739 20791
rect 18739 20757 18748 20791
rect 18696 20748 18748 20757
rect 21824 20791 21876 20800
rect 21824 20757 21833 20791
rect 21833 20757 21867 20791
rect 21867 20757 21876 20791
rect 21824 20748 21876 20757
rect 4266 20646 4318 20698
rect 4330 20646 4382 20698
rect 4394 20646 4446 20698
rect 4458 20646 4510 20698
rect 4522 20646 4574 20698
rect 9579 20646 9631 20698
rect 9643 20646 9695 20698
rect 9707 20646 9759 20698
rect 9771 20646 9823 20698
rect 9835 20646 9887 20698
rect 14892 20646 14944 20698
rect 14956 20646 15008 20698
rect 15020 20646 15072 20698
rect 15084 20646 15136 20698
rect 15148 20646 15200 20698
rect 20205 20646 20257 20698
rect 20269 20646 20321 20698
rect 20333 20646 20385 20698
rect 20397 20646 20449 20698
rect 20461 20646 20513 20698
rect 5448 20544 5500 20596
rect 9956 20544 10008 20596
rect 18236 20544 18288 20596
rect 18696 20544 18748 20596
rect 3976 20408 4028 20460
rect 4804 20204 4856 20256
rect 5356 20451 5408 20460
rect 5356 20417 5365 20451
rect 5365 20417 5399 20451
rect 5399 20417 5408 20451
rect 5356 20408 5408 20417
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 7472 20408 7524 20460
rect 9312 20451 9364 20460
rect 9312 20417 9321 20451
rect 9321 20417 9355 20451
rect 9355 20417 9364 20451
rect 9312 20408 9364 20417
rect 9404 20451 9456 20460
rect 9404 20417 9413 20451
rect 9413 20417 9447 20451
rect 9447 20417 9456 20451
rect 9404 20408 9456 20417
rect 13636 20519 13688 20528
rect 13636 20485 13645 20519
rect 13645 20485 13679 20519
rect 13679 20485 13688 20519
rect 13636 20476 13688 20485
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 15292 20451 15344 20460
rect 15292 20417 15301 20451
rect 15301 20417 15335 20451
rect 15335 20417 15344 20451
rect 15292 20408 15344 20417
rect 17132 20451 17184 20460
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 18328 20408 18380 20460
rect 21824 20408 21876 20460
rect 5632 20340 5684 20392
rect 7196 20383 7248 20392
rect 7196 20349 7205 20383
rect 7205 20349 7239 20383
rect 7239 20349 7248 20383
rect 7196 20340 7248 20349
rect 10784 20340 10836 20392
rect 10968 20383 11020 20392
rect 10968 20349 10977 20383
rect 10977 20349 11011 20383
rect 11011 20349 11020 20383
rect 10968 20340 11020 20349
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 15660 20340 15712 20392
rect 17500 20340 17552 20392
rect 17868 20340 17920 20392
rect 18420 20340 18472 20392
rect 20628 20340 20680 20392
rect 7840 20272 7892 20324
rect 10692 20272 10744 20324
rect 18236 20272 18288 20324
rect 19064 20272 19116 20324
rect 5540 20204 5592 20256
rect 5724 20247 5776 20256
rect 5724 20213 5733 20247
rect 5733 20213 5767 20247
rect 5767 20213 5776 20247
rect 5724 20204 5776 20213
rect 7564 20204 7616 20256
rect 10416 20247 10468 20256
rect 10416 20213 10425 20247
rect 10425 20213 10459 20247
rect 10459 20213 10468 20247
rect 10416 20204 10468 20213
rect 15200 20204 15252 20256
rect 16764 20247 16816 20256
rect 16764 20213 16773 20247
rect 16773 20213 16807 20247
rect 16807 20213 16816 20247
rect 16764 20204 16816 20213
rect 17040 20204 17092 20256
rect 18880 20204 18932 20256
rect 3606 20102 3658 20154
rect 3670 20102 3722 20154
rect 3734 20102 3786 20154
rect 3798 20102 3850 20154
rect 3862 20102 3914 20154
rect 8919 20102 8971 20154
rect 8983 20102 9035 20154
rect 9047 20102 9099 20154
rect 9111 20102 9163 20154
rect 9175 20102 9227 20154
rect 14232 20102 14284 20154
rect 14296 20102 14348 20154
rect 14360 20102 14412 20154
rect 14424 20102 14476 20154
rect 14488 20102 14540 20154
rect 19545 20102 19597 20154
rect 19609 20102 19661 20154
rect 19673 20102 19725 20154
rect 19737 20102 19789 20154
rect 19801 20102 19853 20154
rect 6000 20000 6052 20052
rect 5356 19932 5408 19984
rect 4804 19864 4856 19916
rect 4988 19839 5040 19848
rect 4988 19805 4997 19839
rect 4997 19805 5031 19839
rect 5031 19805 5040 19839
rect 4988 19796 5040 19805
rect 5632 19907 5684 19916
rect 5632 19873 5641 19907
rect 5641 19873 5675 19907
rect 5675 19873 5684 19907
rect 5632 19864 5684 19873
rect 7840 19907 7892 19916
rect 7840 19873 7849 19907
rect 7849 19873 7883 19907
rect 7883 19873 7892 19907
rect 7840 19864 7892 19873
rect 8760 19864 8812 19916
rect 9404 19907 9456 19916
rect 9404 19873 9413 19907
rect 9413 19873 9447 19907
rect 9447 19873 9456 19907
rect 9404 19864 9456 19873
rect 10232 19864 10284 19916
rect 5540 19796 5592 19848
rect 7564 19839 7616 19848
rect 7564 19805 7573 19839
rect 7573 19805 7607 19839
rect 7607 19805 7616 19839
rect 7564 19796 7616 19805
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 10048 19839 10100 19848
rect 10048 19805 10057 19839
rect 10057 19805 10091 19839
rect 10091 19805 10100 19839
rect 13360 20000 13412 20052
rect 15568 20000 15620 20052
rect 13820 19932 13872 19984
rect 12532 19864 12584 19916
rect 13268 19864 13320 19916
rect 13452 19907 13504 19916
rect 13452 19873 13461 19907
rect 13461 19873 13495 19907
rect 13495 19873 13504 19907
rect 13452 19864 13504 19873
rect 17868 20043 17920 20052
rect 17868 20009 17877 20043
rect 17877 20009 17911 20043
rect 17911 20009 17920 20043
rect 17868 20000 17920 20009
rect 18420 19932 18472 19984
rect 10048 19796 10100 19805
rect 7012 19728 7064 19780
rect 10416 19728 10468 19780
rect 12716 19796 12768 19848
rect 14096 19796 14148 19848
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 848 19660 900 19712
rect 7288 19660 7340 19712
rect 11060 19703 11112 19712
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 11244 19660 11296 19712
rect 14464 19771 14516 19780
rect 14464 19737 14473 19771
rect 14473 19737 14507 19771
rect 14507 19737 14516 19771
rect 14464 19728 14516 19737
rect 15476 19728 15528 19780
rect 18328 19907 18380 19916
rect 18328 19873 18337 19907
rect 18337 19873 18371 19907
rect 18371 19873 18380 19907
rect 18328 19864 18380 19873
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 18604 19796 18656 19848
rect 18880 19839 18932 19848
rect 18880 19805 18889 19839
rect 18889 19805 18923 19839
rect 18923 19805 18932 19839
rect 18880 19796 18932 19805
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 13268 19703 13320 19712
rect 13268 19669 13277 19703
rect 13277 19669 13311 19703
rect 13311 19669 13320 19703
rect 13268 19660 13320 19669
rect 14740 19660 14792 19712
rect 17132 19703 17184 19712
rect 17132 19669 17141 19703
rect 17141 19669 17175 19703
rect 17175 19669 17184 19703
rect 17132 19660 17184 19669
rect 18512 19703 18564 19712
rect 18512 19669 18521 19703
rect 18521 19669 18555 19703
rect 18555 19669 18564 19703
rect 18512 19660 18564 19669
rect 21824 19703 21876 19712
rect 21824 19669 21833 19703
rect 21833 19669 21867 19703
rect 21867 19669 21876 19703
rect 21824 19660 21876 19669
rect 4266 19558 4318 19610
rect 4330 19558 4382 19610
rect 4394 19558 4446 19610
rect 4458 19558 4510 19610
rect 4522 19558 4574 19610
rect 9579 19558 9631 19610
rect 9643 19558 9695 19610
rect 9707 19558 9759 19610
rect 9771 19558 9823 19610
rect 9835 19558 9887 19610
rect 14892 19558 14944 19610
rect 14956 19558 15008 19610
rect 15020 19558 15072 19610
rect 15084 19558 15136 19610
rect 15148 19558 15200 19610
rect 20205 19558 20257 19610
rect 20269 19558 20321 19610
rect 20333 19558 20385 19610
rect 20397 19558 20449 19610
rect 20461 19558 20513 19610
rect 7288 19499 7340 19508
rect 7288 19465 7297 19499
rect 7297 19465 7331 19499
rect 7331 19465 7340 19499
rect 7288 19456 7340 19465
rect 7380 19499 7432 19508
rect 7380 19465 7389 19499
rect 7389 19465 7423 19499
rect 7423 19465 7432 19499
rect 7380 19456 7432 19465
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 10140 19499 10192 19508
rect 10140 19465 10149 19499
rect 10149 19465 10183 19499
rect 10183 19465 10192 19499
rect 10140 19456 10192 19465
rect 7472 19388 7524 19440
rect 10784 19431 10836 19440
rect 10784 19397 10793 19431
rect 10793 19397 10827 19431
rect 10827 19397 10836 19431
rect 10784 19388 10836 19397
rect 11152 19456 11204 19508
rect 12808 19456 12860 19508
rect 13820 19456 13872 19508
rect 14004 19499 14056 19508
rect 14004 19465 14013 19499
rect 14013 19465 14047 19499
rect 14047 19465 14056 19499
rect 14004 19456 14056 19465
rect 11244 19388 11296 19440
rect 4988 19320 5040 19372
rect 2872 19252 2924 19304
rect 4160 19252 4212 19304
rect 4804 19252 4856 19304
rect 5816 19184 5868 19236
rect 8576 19320 8628 19372
rect 7840 19184 7892 19236
rect 10048 19252 10100 19304
rect 11060 19320 11112 19372
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 13544 19320 13596 19372
rect 13912 19320 13964 19372
rect 14648 19499 14700 19508
rect 14648 19465 14657 19499
rect 14657 19465 14691 19499
rect 14691 19465 14700 19499
rect 14648 19456 14700 19465
rect 14740 19499 14792 19508
rect 14740 19465 14749 19499
rect 14749 19465 14783 19499
rect 14783 19465 14792 19499
rect 14740 19456 14792 19465
rect 15844 19456 15896 19508
rect 17040 19499 17092 19508
rect 17040 19465 17049 19499
rect 17049 19465 17083 19499
rect 17083 19465 17092 19499
rect 17040 19456 17092 19465
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 21640 19456 21692 19508
rect 22008 19363 22060 19372
rect 22008 19329 22017 19363
rect 22017 19329 22051 19363
rect 22051 19329 22060 19363
rect 22008 19320 22060 19329
rect 13176 19295 13228 19304
rect 13176 19261 13185 19295
rect 13185 19261 13219 19295
rect 13219 19261 13228 19295
rect 13176 19252 13228 19261
rect 13268 19252 13320 19304
rect 14464 19252 14516 19304
rect 17408 19252 17460 19304
rect 10232 19184 10284 19236
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 5908 19116 5960 19168
rect 7380 19116 7432 19168
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8392 19116 8444 19125
rect 9772 19159 9824 19168
rect 9772 19125 9781 19159
rect 9781 19125 9815 19159
rect 9815 19125 9824 19159
rect 9772 19116 9824 19125
rect 10968 19159 11020 19168
rect 10968 19125 10977 19159
rect 10977 19125 11011 19159
rect 11011 19125 11020 19159
rect 10968 19116 11020 19125
rect 3606 19014 3658 19066
rect 3670 19014 3722 19066
rect 3734 19014 3786 19066
rect 3798 19014 3850 19066
rect 3862 19014 3914 19066
rect 8919 19014 8971 19066
rect 8983 19014 9035 19066
rect 9047 19014 9099 19066
rect 9111 19014 9163 19066
rect 9175 19014 9227 19066
rect 14232 19014 14284 19066
rect 14296 19014 14348 19066
rect 14360 19014 14412 19066
rect 14424 19014 14476 19066
rect 14488 19014 14540 19066
rect 19545 19014 19597 19066
rect 19609 19014 19661 19066
rect 19673 19014 19725 19066
rect 19737 19014 19789 19066
rect 19801 19014 19853 19066
rect 4988 18912 5040 18964
rect 848 18708 900 18760
rect 2504 18776 2556 18828
rect 7840 18912 7892 18964
rect 10140 18912 10192 18964
rect 6644 18844 6696 18896
rect 14096 18844 14148 18896
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 8576 18819 8628 18828
rect 8576 18785 8585 18819
rect 8585 18785 8619 18819
rect 8619 18785 8628 18819
rect 8576 18776 8628 18785
rect 2964 18708 3016 18760
rect 5172 18751 5224 18760
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 5908 18751 5960 18760
rect 5908 18717 5917 18751
rect 5917 18717 5951 18751
rect 5951 18717 5960 18751
rect 5908 18708 5960 18717
rect 9772 18708 9824 18760
rect 4804 18640 4856 18692
rect 6552 18683 6604 18692
rect 6552 18649 6561 18683
rect 6561 18649 6595 18683
rect 6595 18649 6604 18683
rect 6552 18640 6604 18649
rect 10416 18819 10468 18828
rect 10416 18785 10425 18819
rect 10425 18785 10459 18819
rect 10459 18785 10468 18819
rect 10416 18776 10468 18785
rect 10232 18751 10284 18760
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 18144 18751 18196 18760
rect 18144 18717 18153 18751
rect 18153 18717 18187 18751
rect 18187 18717 18196 18751
rect 18144 18708 18196 18717
rect 22008 18751 22060 18760
rect 22008 18717 22017 18751
rect 22017 18717 22051 18751
rect 22051 18717 22060 18751
rect 22008 18708 22060 18717
rect 12532 18640 12584 18692
rect 1860 18572 1912 18624
rect 2780 18615 2832 18624
rect 2780 18581 2789 18615
rect 2789 18581 2823 18615
rect 2823 18581 2832 18615
rect 2780 18572 2832 18581
rect 3332 18572 3384 18624
rect 5632 18572 5684 18624
rect 7564 18572 7616 18624
rect 20996 18572 21048 18624
rect 4266 18470 4318 18522
rect 4330 18470 4382 18522
rect 4394 18470 4446 18522
rect 4458 18470 4510 18522
rect 4522 18470 4574 18522
rect 9579 18470 9631 18522
rect 9643 18470 9695 18522
rect 9707 18470 9759 18522
rect 9771 18470 9823 18522
rect 9835 18470 9887 18522
rect 14892 18470 14944 18522
rect 14956 18470 15008 18522
rect 15020 18470 15072 18522
rect 15084 18470 15136 18522
rect 15148 18470 15200 18522
rect 20205 18470 20257 18522
rect 20269 18470 20321 18522
rect 20333 18470 20385 18522
rect 20397 18470 20449 18522
rect 20461 18470 20513 18522
rect 1584 18368 1636 18420
rect 2596 18368 2648 18420
rect 2780 18368 2832 18420
rect 3332 18411 3384 18420
rect 3332 18377 3341 18411
rect 3341 18377 3375 18411
rect 3375 18377 3384 18411
rect 3332 18368 3384 18377
rect 4804 18300 4856 18352
rect 5632 18411 5684 18420
rect 5632 18377 5641 18411
rect 5641 18377 5675 18411
rect 5675 18377 5684 18411
rect 5632 18368 5684 18377
rect 5724 18411 5776 18420
rect 5724 18377 5733 18411
rect 5733 18377 5767 18411
rect 5767 18377 5776 18411
rect 5724 18368 5776 18377
rect 7196 18411 7248 18420
rect 7196 18377 7205 18411
rect 7205 18377 7239 18411
rect 7239 18377 7248 18411
rect 7196 18368 7248 18377
rect 7932 18368 7984 18420
rect 13544 18411 13596 18420
rect 13544 18377 13553 18411
rect 13553 18377 13587 18411
rect 13587 18377 13596 18411
rect 13544 18368 13596 18377
rect 16672 18368 16724 18420
rect 18144 18411 18196 18420
rect 18144 18377 18153 18411
rect 18153 18377 18187 18411
rect 18187 18377 18196 18411
rect 18144 18368 18196 18377
rect 6920 18300 6972 18352
rect 13820 18300 13872 18352
rect 14096 18300 14148 18352
rect 17040 18300 17092 18352
rect 19340 18300 19392 18352
rect 19432 18300 19484 18352
rect 19892 18343 19944 18352
rect 19892 18309 19901 18343
rect 19901 18309 19935 18343
rect 19935 18309 19944 18343
rect 19892 18300 19944 18309
rect 1860 18275 1912 18284
rect 1860 18241 1904 18275
rect 1904 18241 1912 18275
rect 1860 18232 1912 18241
rect 2412 18207 2464 18216
rect 2412 18173 2421 18207
rect 2421 18173 2455 18207
rect 2455 18173 2464 18207
rect 2412 18164 2464 18173
rect 2872 18232 2924 18284
rect 4068 18232 4120 18284
rect 4896 18275 4948 18284
rect 4896 18241 4905 18275
rect 4905 18241 4939 18275
rect 4939 18241 4948 18275
rect 4896 18232 4948 18241
rect 5724 18232 5776 18284
rect 6644 18232 6696 18284
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 7564 18275 7616 18284
rect 7564 18241 7573 18275
rect 7573 18241 7607 18275
rect 7607 18241 7616 18275
rect 7564 18232 7616 18241
rect 13360 18275 13412 18284
rect 13360 18241 13369 18275
rect 13369 18241 13403 18275
rect 13403 18241 13412 18275
rect 13360 18232 13412 18241
rect 13636 18275 13688 18284
rect 13636 18241 13645 18275
rect 13645 18241 13679 18275
rect 13679 18241 13688 18275
rect 13636 18232 13688 18241
rect 13912 18275 13964 18284
rect 13912 18241 13921 18275
rect 13921 18241 13955 18275
rect 13955 18241 13964 18275
rect 13912 18232 13964 18241
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 2964 18096 3016 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 1952 18028 2004 18080
rect 3976 18164 4028 18216
rect 5816 18164 5868 18216
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 6000 18096 6052 18148
rect 12716 18139 12768 18148
rect 12716 18105 12725 18139
rect 12725 18105 12759 18139
rect 12759 18105 12768 18139
rect 12716 18096 12768 18105
rect 13268 18096 13320 18148
rect 18052 18275 18104 18284
rect 18052 18241 18061 18275
rect 18061 18241 18095 18275
rect 18095 18241 18104 18275
rect 18052 18232 18104 18241
rect 20996 18275 21048 18284
rect 20996 18241 21004 18275
rect 21004 18241 21048 18275
rect 20996 18232 21048 18241
rect 21088 18232 21140 18284
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 18420 18164 18472 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 4160 18028 4212 18080
rect 4896 18028 4948 18080
rect 6184 18028 6236 18080
rect 17316 18096 17368 18148
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 3606 17926 3658 17978
rect 3670 17926 3722 17978
rect 3734 17926 3786 17978
rect 3798 17926 3850 17978
rect 3862 17926 3914 17978
rect 8919 17926 8971 17978
rect 8983 17926 9035 17978
rect 9047 17926 9099 17978
rect 9111 17926 9163 17978
rect 9175 17926 9227 17978
rect 14232 17926 14284 17978
rect 14296 17926 14348 17978
rect 14360 17926 14412 17978
rect 14424 17926 14476 17978
rect 14488 17926 14540 17978
rect 19545 17926 19597 17978
rect 19609 17926 19661 17978
rect 19673 17926 19725 17978
rect 19737 17926 19789 17978
rect 19801 17926 19853 17978
rect 2412 17824 2464 17876
rect 4712 17824 4764 17876
rect 6920 17867 6972 17876
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 7380 17824 7432 17876
rect 13360 17824 13412 17876
rect 18052 17867 18104 17876
rect 18052 17833 18061 17867
rect 18061 17833 18095 17867
rect 18095 17833 18104 17867
rect 18052 17824 18104 17833
rect 2964 17756 3016 17808
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 1952 17731 2004 17740
rect 1952 17697 1961 17731
rect 1961 17697 1995 17731
rect 1995 17697 2004 17731
rect 1952 17688 2004 17697
rect 4068 17756 4120 17808
rect 1860 17620 1912 17672
rect 2596 17663 2648 17672
rect 2596 17629 2630 17663
rect 2630 17629 2648 17663
rect 2596 17620 2648 17629
rect 3976 17620 4028 17672
rect 4896 17731 4948 17740
rect 4896 17697 4905 17731
rect 4905 17697 4939 17731
rect 4939 17697 4948 17731
rect 4896 17688 4948 17697
rect 5172 17688 5224 17740
rect 5816 17731 5868 17740
rect 5816 17697 5825 17731
rect 5825 17697 5859 17731
rect 5859 17697 5868 17731
rect 5816 17688 5868 17697
rect 8852 17688 8904 17740
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 6000 17663 6052 17672
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 2504 17484 2556 17536
rect 7564 17620 7616 17672
rect 8944 17663 8996 17672
rect 8944 17629 8953 17663
rect 8953 17629 8987 17663
rect 8987 17629 8996 17663
rect 8944 17620 8996 17629
rect 10968 17688 11020 17740
rect 7748 17552 7800 17604
rect 10140 17552 10192 17604
rect 11152 17595 11204 17604
rect 11152 17561 11161 17595
rect 11161 17561 11195 17595
rect 11195 17561 11204 17595
rect 11152 17552 11204 17561
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 13452 17756 13504 17808
rect 12716 17620 12768 17672
rect 16396 17688 16448 17740
rect 18604 17688 18656 17740
rect 19524 17731 19576 17740
rect 19524 17697 19533 17731
rect 19533 17697 19567 17731
rect 19567 17697 19576 17731
rect 19524 17688 19576 17697
rect 20628 17688 20680 17740
rect 18512 17620 18564 17672
rect 19892 17620 19944 17672
rect 21824 17620 21876 17672
rect 18788 17552 18840 17604
rect 19064 17595 19116 17604
rect 19064 17561 19073 17595
rect 19073 17561 19107 17595
rect 19107 17561 19116 17595
rect 19064 17552 19116 17561
rect 8668 17484 8720 17536
rect 15292 17484 15344 17536
rect 18696 17527 18748 17536
rect 18696 17493 18705 17527
rect 18705 17493 18739 17527
rect 18739 17493 18748 17527
rect 18696 17484 18748 17493
rect 4266 17382 4318 17434
rect 4330 17382 4382 17434
rect 4394 17382 4446 17434
rect 4458 17382 4510 17434
rect 4522 17382 4574 17434
rect 9579 17382 9631 17434
rect 9643 17382 9695 17434
rect 9707 17382 9759 17434
rect 9771 17382 9823 17434
rect 9835 17382 9887 17434
rect 14892 17382 14944 17434
rect 14956 17382 15008 17434
rect 15020 17382 15072 17434
rect 15084 17382 15136 17434
rect 15148 17382 15200 17434
rect 20205 17382 20257 17434
rect 20269 17382 20321 17434
rect 20333 17382 20385 17434
rect 20397 17382 20449 17434
rect 20461 17382 20513 17434
rect 8852 17323 8904 17332
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 8944 17323 8996 17332
rect 8944 17289 8953 17323
rect 8953 17289 8987 17323
rect 8987 17289 8996 17323
rect 8944 17280 8996 17289
rect 11152 17280 11204 17332
rect 10508 17212 10560 17264
rect 6184 17187 6236 17196
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 12716 17212 12768 17264
rect 12900 17212 12952 17264
rect 15292 17280 15344 17332
rect 8484 17076 8536 17128
rect 10140 17076 10192 17128
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 848 17008 900 17060
rect 17960 17280 18012 17332
rect 18788 17323 18840 17332
rect 18788 17289 18797 17323
rect 18797 17289 18831 17323
rect 18831 17289 18840 17323
rect 18788 17280 18840 17289
rect 19064 17280 19116 17332
rect 19340 17323 19392 17332
rect 19340 17289 19349 17323
rect 19349 17289 19383 17323
rect 19383 17289 19392 17323
rect 19340 17280 19392 17289
rect 15752 17144 15804 17196
rect 18604 17187 18656 17196
rect 18604 17153 18613 17187
rect 18613 17153 18647 17187
rect 18647 17153 18656 17187
rect 18604 17144 18656 17153
rect 19524 17187 19576 17196
rect 19524 17153 19533 17187
rect 19533 17153 19567 17187
rect 19567 17153 19576 17187
rect 19524 17144 19576 17153
rect 21364 17187 21416 17196
rect 21364 17153 21373 17187
rect 21373 17153 21407 17187
rect 21407 17153 21416 17187
rect 21364 17144 21416 17153
rect 12992 17076 13044 17128
rect 13544 17076 13596 17128
rect 13728 17076 13780 17128
rect 10784 17008 10836 17060
rect 12532 17008 12584 17060
rect 18512 17076 18564 17128
rect 19892 17076 19944 17128
rect 21548 17051 21600 17060
rect 21548 17017 21557 17051
rect 21557 17017 21591 17051
rect 21591 17017 21600 17051
rect 21548 17008 21600 17017
rect 8300 16940 8352 16992
rect 3606 16838 3658 16890
rect 3670 16838 3722 16890
rect 3734 16838 3786 16890
rect 3798 16838 3850 16890
rect 3862 16838 3914 16890
rect 8919 16838 8971 16890
rect 8983 16838 9035 16890
rect 9047 16838 9099 16890
rect 9111 16838 9163 16890
rect 9175 16838 9227 16890
rect 14232 16838 14284 16890
rect 14296 16838 14348 16890
rect 14360 16838 14412 16890
rect 14424 16838 14476 16890
rect 14488 16838 14540 16890
rect 19545 16838 19597 16890
rect 19609 16838 19661 16890
rect 19673 16838 19725 16890
rect 19737 16838 19789 16890
rect 19801 16838 19853 16890
rect 10692 16736 10744 16788
rect 8484 16668 8536 16720
rect 8300 16643 8352 16652
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 8576 16600 8628 16652
rect 848 16532 900 16584
rect 5632 16575 5684 16584
rect 5632 16541 5641 16575
rect 5641 16541 5675 16575
rect 5675 16541 5684 16575
rect 5632 16532 5684 16541
rect 6736 16464 6788 16516
rect 7748 16575 7800 16584
rect 7748 16541 7757 16575
rect 7757 16541 7791 16575
rect 7791 16541 7800 16575
rect 7748 16532 7800 16541
rect 10508 16643 10560 16652
rect 10508 16609 10517 16643
rect 10517 16609 10551 16643
rect 10551 16609 10560 16643
rect 10508 16600 10560 16609
rect 12992 16779 13044 16788
rect 12992 16745 13001 16779
rect 13001 16745 13035 16779
rect 13035 16745 13044 16779
rect 12992 16736 13044 16745
rect 15844 16736 15896 16788
rect 12900 16668 12952 16720
rect 12624 16600 12676 16652
rect 13176 16600 13228 16652
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 15292 16532 15344 16584
rect 16304 16575 16356 16584
rect 16304 16541 16313 16575
rect 16313 16541 16347 16575
rect 16347 16541 16356 16575
rect 16304 16532 16356 16541
rect 21088 16532 21140 16584
rect 22008 16575 22060 16584
rect 22008 16541 22017 16575
rect 22017 16541 22051 16575
rect 22051 16541 22060 16575
rect 22008 16532 22060 16541
rect 2044 16396 2096 16448
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 7472 16396 7524 16448
rect 10784 16507 10836 16516
rect 10784 16473 10793 16507
rect 10793 16473 10827 16507
rect 10827 16473 10836 16507
rect 10784 16464 10836 16473
rect 10508 16396 10560 16448
rect 13820 16464 13872 16516
rect 15384 16507 15436 16516
rect 15384 16473 15393 16507
rect 15393 16473 15427 16507
rect 15427 16473 15436 16507
rect 15384 16464 15436 16473
rect 12532 16439 12584 16448
rect 12532 16405 12541 16439
rect 12541 16405 12575 16439
rect 12575 16405 12584 16439
rect 12532 16396 12584 16405
rect 13544 16439 13596 16448
rect 13544 16405 13553 16439
rect 13553 16405 13587 16439
rect 13587 16405 13596 16439
rect 13544 16396 13596 16405
rect 15568 16396 15620 16448
rect 21364 16464 21416 16516
rect 21732 16396 21784 16448
rect 4266 16294 4318 16346
rect 4330 16294 4382 16346
rect 4394 16294 4446 16346
rect 4458 16294 4510 16346
rect 4522 16294 4574 16346
rect 9579 16294 9631 16346
rect 9643 16294 9695 16346
rect 9707 16294 9759 16346
rect 9771 16294 9823 16346
rect 9835 16294 9887 16346
rect 14892 16294 14944 16346
rect 14956 16294 15008 16346
rect 15020 16294 15072 16346
rect 15084 16294 15136 16346
rect 15148 16294 15200 16346
rect 20205 16294 20257 16346
rect 20269 16294 20321 16346
rect 20333 16294 20385 16346
rect 20397 16294 20449 16346
rect 20461 16294 20513 16346
rect 3976 16235 4028 16244
rect 3976 16201 3985 16235
rect 3985 16201 4019 16235
rect 4019 16201 4028 16235
rect 3976 16192 4028 16201
rect 5632 16192 5684 16244
rect 6828 16235 6880 16244
rect 6828 16201 6837 16235
rect 6837 16201 6871 16235
rect 6871 16201 6880 16235
rect 6828 16192 6880 16201
rect 10508 16192 10560 16244
rect 12532 16192 12584 16244
rect 13544 16192 13596 16244
rect 15384 16192 15436 16244
rect 16304 16192 16356 16244
rect 2412 16099 2464 16108
rect 2412 16065 2421 16099
rect 2421 16065 2455 16099
rect 2455 16065 2464 16099
rect 2412 16056 2464 16065
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 6276 16124 6328 16176
rect 6736 16167 6788 16176
rect 6736 16133 6745 16167
rect 6745 16133 6779 16167
rect 6779 16133 6788 16167
rect 6736 16124 6788 16133
rect 3424 16056 3476 16108
rect 4620 16056 4672 16108
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 5632 16056 5684 16065
rect 2872 15988 2924 16040
rect 3976 15988 4028 16040
rect 4160 15988 4212 16040
rect 5356 15988 5408 16040
rect 6460 15988 6512 16040
rect 6092 15920 6144 15972
rect 6184 15920 6236 15972
rect 848 15852 900 15904
rect 4068 15852 4120 15904
rect 5448 15852 5500 15904
rect 5908 15852 5960 15904
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 10876 16056 10928 16108
rect 11704 16099 11756 16108
rect 11704 16065 11712 16099
rect 11712 16065 11756 16099
rect 11704 16056 11756 16065
rect 13820 16124 13872 16176
rect 14556 16124 14608 16176
rect 13452 16099 13504 16108
rect 13452 16065 13486 16099
rect 13486 16065 13504 16099
rect 13452 16056 13504 16065
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 18328 16056 18380 16108
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 10600 15988 10652 16040
rect 12624 15988 12676 16040
rect 15752 16031 15804 16040
rect 15752 15997 15761 16031
rect 15761 15997 15795 16031
rect 15795 15997 15804 16031
rect 15752 15988 15804 15997
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 17408 15988 17460 16040
rect 12164 15920 12216 15972
rect 16304 15920 16356 15972
rect 18880 15920 18932 15972
rect 7472 15852 7524 15904
rect 10508 15852 10560 15904
rect 16212 15895 16264 15904
rect 16212 15861 16221 15895
rect 16221 15861 16255 15895
rect 16255 15861 16264 15895
rect 16212 15852 16264 15861
rect 21088 15852 21140 15904
rect 3606 15750 3658 15802
rect 3670 15750 3722 15802
rect 3734 15750 3786 15802
rect 3798 15750 3850 15802
rect 3862 15750 3914 15802
rect 8919 15750 8971 15802
rect 8983 15750 9035 15802
rect 9047 15750 9099 15802
rect 9111 15750 9163 15802
rect 9175 15750 9227 15802
rect 14232 15750 14284 15802
rect 14296 15750 14348 15802
rect 14360 15750 14412 15802
rect 14424 15750 14476 15802
rect 14488 15750 14540 15802
rect 19545 15750 19597 15802
rect 19609 15750 19661 15802
rect 19673 15750 19725 15802
rect 19737 15750 19789 15802
rect 19801 15750 19853 15802
rect 2412 15691 2464 15700
rect 2412 15657 2421 15691
rect 2421 15657 2455 15691
rect 2455 15657 2464 15691
rect 2412 15648 2464 15657
rect 2596 15648 2648 15700
rect 5908 15691 5960 15700
rect 5908 15657 5917 15691
rect 5917 15657 5951 15691
rect 5951 15657 5960 15691
rect 5908 15648 5960 15657
rect 6092 15648 6144 15700
rect 7748 15691 7800 15700
rect 7748 15657 7757 15691
rect 7757 15657 7791 15691
rect 7791 15657 7800 15691
rect 7748 15648 7800 15657
rect 10784 15648 10836 15700
rect 11888 15648 11940 15700
rect 15752 15691 15804 15700
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 18420 15691 18472 15700
rect 18420 15657 18429 15691
rect 18429 15657 18463 15691
rect 18463 15657 18472 15691
rect 18420 15648 18472 15657
rect 19340 15648 19392 15700
rect 2872 15580 2924 15632
rect 1768 15512 1820 15564
rect 2136 15512 2188 15564
rect 4160 15580 4212 15632
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 5816 15580 5868 15632
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 8576 15580 8628 15632
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 3976 15444 4028 15496
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 2044 15419 2096 15428
rect 2044 15385 2053 15419
rect 2053 15385 2087 15419
rect 2087 15385 2096 15419
rect 2044 15376 2096 15385
rect 1952 15351 2004 15360
rect 1952 15317 1961 15351
rect 1961 15317 1995 15351
rect 1995 15317 2004 15351
rect 1952 15308 2004 15317
rect 2136 15308 2188 15360
rect 2872 15308 2924 15360
rect 4160 15351 4212 15360
rect 4160 15317 4169 15351
rect 4169 15317 4203 15351
rect 4203 15317 4212 15351
rect 4160 15308 4212 15317
rect 7748 15376 7800 15428
rect 10508 15512 10560 15564
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 10876 15487 10928 15496
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 16304 15555 16356 15564
rect 16304 15521 16313 15555
rect 16313 15521 16347 15555
rect 16347 15521 16356 15555
rect 16304 15512 16356 15521
rect 19156 15512 19208 15564
rect 8484 15308 8536 15360
rect 10508 15376 10560 15428
rect 10692 15376 10744 15428
rect 13636 15444 13688 15496
rect 18788 15487 18840 15496
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 21088 15444 21140 15496
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 10600 15308 10652 15360
rect 16120 15351 16172 15360
rect 16120 15317 16129 15351
rect 16129 15317 16163 15351
rect 16163 15317 16172 15351
rect 16120 15308 16172 15317
rect 21180 15308 21232 15360
rect 21824 15351 21876 15360
rect 21824 15317 21833 15351
rect 21833 15317 21867 15351
rect 21867 15317 21876 15351
rect 21824 15308 21876 15317
rect 4266 15206 4318 15258
rect 4330 15206 4382 15258
rect 4394 15206 4446 15258
rect 4458 15206 4510 15258
rect 4522 15206 4574 15258
rect 9579 15206 9631 15258
rect 9643 15206 9695 15258
rect 9707 15206 9759 15258
rect 9771 15206 9823 15258
rect 9835 15206 9887 15258
rect 14892 15206 14944 15258
rect 14956 15206 15008 15258
rect 15020 15206 15072 15258
rect 15084 15206 15136 15258
rect 15148 15206 15200 15258
rect 20205 15206 20257 15258
rect 20269 15206 20321 15258
rect 20333 15206 20385 15258
rect 20397 15206 20449 15258
rect 20461 15206 20513 15258
rect 1952 15104 2004 15156
rect 3424 15104 3476 15156
rect 4160 15104 4212 15156
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 8576 15104 8628 15156
rect 13636 15104 13688 15156
rect 18328 15147 18380 15156
rect 18328 15113 18337 15147
rect 18337 15113 18371 15147
rect 18371 15113 18380 15147
rect 18328 15104 18380 15113
rect 2044 15011 2096 15020
rect 2044 14977 2062 15011
rect 2062 14977 2096 15011
rect 2044 14968 2096 14977
rect 2412 14900 2464 14952
rect 2596 14968 2648 15020
rect 4620 15036 4672 15088
rect 4712 14900 4764 14952
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 8116 15011 8168 15020
rect 8116 14977 8125 15011
rect 8125 14977 8159 15011
rect 8159 14977 8168 15011
rect 8116 14968 8168 14977
rect 9404 14968 9456 15020
rect 5632 14943 5684 14952
rect 5632 14909 5641 14943
rect 5641 14909 5675 14943
rect 5675 14909 5684 14943
rect 5632 14900 5684 14909
rect 8300 14943 8352 14952
rect 8300 14909 8309 14943
rect 8309 14909 8343 14943
rect 8343 14909 8352 14943
rect 8300 14900 8352 14909
rect 8484 14832 8536 14884
rect 8760 14900 8812 14952
rect 15844 15036 15896 15088
rect 12992 14968 13044 15020
rect 16488 14968 16540 15020
rect 13084 14900 13136 14952
rect 15476 14900 15528 14952
rect 16120 14900 16172 14952
rect 19432 15036 19484 15088
rect 21088 15147 21140 15156
rect 21088 15113 21097 15147
rect 21097 15113 21131 15147
rect 21131 15113 21140 15147
rect 21088 15104 21140 15113
rect 21180 15147 21232 15156
rect 21180 15113 21189 15147
rect 21189 15113 21223 15147
rect 21223 15113 21232 15147
rect 21180 15104 21232 15113
rect 19248 14968 19300 15020
rect 20720 15036 20772 15088
rect 21824 15036 21876 15088
rect 20076 14968 20128 15020
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 19156 14943 19208 14952
rect 19156 14909 19165 14943
rect 19165 14909 19199 14943
rect 19199 14909 19208 14943
rect 19156 14900 19208 14909
rect 20352 14943 20404 14952
rect 20352 14909 20361 14943
rect 20361 14909 20395 14943
rect 20395 14909 20404 14943
rect 20352 14900 20404 14909
rect 20536 14968 20588 15020
rect 20628 14900 20680 14952
rect 19892 14832 19944 14884
rect 12900 14764 12952 14816
rect 13544 14764 13596 14816
rect 3606 14662 3658 14714
rect 3670 14662 3722 14714
rect 3734 14662 3786 14714
rect 3798 14662 3850 14714
rect 3862 14662 3914 14714
rect 8919 14662 8971 14714
rect 8983 14662 9035 14714
rect 9047 14662 9099 14714
rect 9111 14662 9163 14714
rect 9175 14662 9227 14714
rect 14232 14662 14284 14714
rect 14296 14662 14348 14714
rect 14360 14662 14412 14714
rect 14424 14662 14476 14714
rect 14488 14662 14540 14714
rect 19545 14662 19597 14714
rect 19609 14662 19661 14714
rect 19673 14662 19725 14714
rect 19737 14662 19789 14714
rect 19801 14662 19853 14714
rect 6460 14560 6512 14612
rect 8760 14560 8812 14612
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 9496 14560 9548 14612
rect 1676 14492 1728 14544
rect 9680 14492 9732 14544
rect 10140 14603 10192 14612
rect 10140 14569 10149 14603
rect 10149 14569 10183 14603
rect 10183 14569 10192 14603
rect 10140 14560 10192 14569
rect 13084 14603 13136 14612
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 9864 14492 9916 14544
rect 10232 14492 10284 14544
rect 5816 14424 5868 14476
rect 848 14356 900 14408
rect 5356 14356 5408 14408
rect 8300 14424 8352 14476
rect 6092 14356 6144 14408
rect 6552 14356 6604 14408
rect 9220 14356 9272 14408
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 5724 14263 5776 14272
rect 5724 14229 5733 14263
rect 5733 14229 5767 14263
rect 5767 14229 5776 14263
rect 5724 14220 5776 14229
rect 9496 14288 9548 14340
rect 6368 14220 6420 14272
rect 8668 14220 8720 14272
rect 9404 14220 9456 14272
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 13728 14467 13780 14476
rect 13728 14433 13737 14467
rect 13737 14433 13771 14467
rect 13771 14433 13780 14467
rect 13728 14424 13780 14433
rect 12440 14356 12492 14408
rect 15384 14560 15436 14612
rect 15476 14603 15528 14612
rect 15476 14569 15485 14603
rect 15485 14569 15519 14603
rect 15519 14569 15528 14603
rect 15476 14560 15528 14569
rect 15660 14560 15712 14612
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 15292 14492 15344 14544
rect 16028 14492 16080 14544
rect 16304 14560 16356 14612
rect 16488 14603 16540 14612
rect 16488 14569 16497 14603
rect 16497 14569 16531 14603
rect 16531 14569 16540 14603
rect 16488 14560 16540 14569
rect 19248 14603 19300 14612
rect 19248 14569 19257 14603
rect 19257 14569 19291 14603
rect 19291 14569 19300 14603
rect 19248 14560 19300 14569
rect 20352 14560 20404 14612
rect 13360 14220 13412 14272
rect 13728 14220 13780 14272
rect 19432 14492 19484 14544
rect 16304 14424 16356 14476
rect 17316 14356 17368 14408
rect 19340 14356 19392 14408
rect 19892 14356 19944 14408
rect 20720 14356 20772 14408
rect 22008 14399 22060 14408
rect 22008 14365 22017 14399
rect 22017 14365 22051 14399
rect 22051 14365 22060 14399
rect 22008 14356 22060 14365
rect 15384 14220 15436 14272
rect 16672 14220 16724 14272
rect 18880 14331 18932 14340
rect 18880 14297 18889 14331
rect 18889 14297 18923 14331
rect 18923 14297 18932 14331
rect 18880 14288 18932 14297
rect 17316 14220 17368 14272
rect 20536 14220 20588 14272
rect 4266 14118 4318 14170
rect 4330 14118 4382 14170
rect 4394 14118 4446 14170
rect 4458 14118 4510 14170
rect 4522 14118 4574 14170
rect 9579 14118 9631 14170
rect 9643 14118 9695 14170
rect 9707 14118 9759 14170
rect 9771 14118 9823 14170
rect 9835 14118 9887 14170
rect 14892 14118 14944 14170
rect 14956 14118 15008 14170
rect 15020 14118 15072 14170
rect 15084 14118 15136 14170
rect 15148 14118 15200 14170
rect 20205 14118 20257 14170
rect 20269 14118 20321 14170
rect 20333 14118 20385 14170
rect 20397 14118 20449 14170
rect 20461 14118 20513 14170
rect 1584 14016 1636 14068
rect 9312 14016 9364 14068
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 12992 14059 13044 14068
rect 12992 14025 13001 14059
rect 13001 14025 13035 14059
rect 13035 14025 13044 14059
rect 12992 14016 13044 14025
rect 14648 14016 14700 14068
rect 16672 14059 16724 14068
rect 16672 14025 16681 14059
rect 16681 14025 16715 14059
rect 16715 14025 16724 14059
rect 16672 14016 16724 14025
rect 10048 13948 10100 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 4712 13880 4764 13932
rect 4896 13880 4948 13932
rect 5264 13880 5316 13932
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 5908 13923 5960 13932
rect 5908 13889 5917 13923
rect 5917 13889 5951 13923
rect 5951 13889 5960 13923
rect 5908 13880 5960 13889
rect 8208 13880 8260 13932
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 9680 13880 9732 13932
rect 11520 13948 11572 14000
rect 12348 13948 12400 14000
rect 1676 13812 1728 13864
rect 6092 13812 6144 13864
rect 6368 13855 6420 13864
rect 6368 13821 6377 13855
rect 6377 13821 6411 13855
rect 6411 13821 6420 13855
rect 6368 13812 6420 13821
rect 5908 13744 5960 13796
rect 8116 13812 8168 13864
rect 9312 13812 9364 13864
rect 9956 13812 10008 13864
rect 10600 13812 10652 13864
rect 10048 13744 10100 13796
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 15292 13812 15344 13864
rect 15476 13812 15528 13864
rect 17316 14016 17368 14068
rect 18880 14016 18932 14068
rect 21640 13948 21692 14000
rect 19892 13880 19944 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 17132 13744 17184 13796
rect 19432 13812 19484 13864
rect 20628 13744 20680 13796
rect 10324 13676 10376 13728
rect 21824 13719 21876 13728
rect 21824 13685 21833 13719
rect 21833 13685 21867 13719
rect 21867 13685 21876 13719
rect 21824 13676 21876 13685
rect 3606 13574 3658 13626
rect 3670 13574 3722 13626
rect 3734 13574 3786 13626
rect 3798 13574 3850 13626
rect 3862 13574 3914 13626
rect 8919 13574 8971 13626
rect 8983 13574 9035 13626
rect 9047 13574 9099 13626
rect 9111 13574 9163 13626
rect 9175 13574 9227 13626
rect 14232 13574 14284 13626
rect 14296 13574 14348 13626
rect 14360 13574 14412 13626
rect 14424 13574 14476 13626
rect 14488 13574 14540 13626
rect 19545 13574 19597 13626
rect 19609 13574 19661 13626
rect 19673 13574 19725 13626
rect 19737 13574 19789 13626
rect 19801 13574 19853 13626
rect 5356 13472 5408 13524
rect 5724 13472 5776 13524
rect 8208 13472 8260 13524
rect 12624 13472 12676 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 5908 13404 5960 13456
rect 9680 13404 9732 13456
rect 848 13268 900 13320
rect 5080 13336 5132 13388
rect 6000 13379 6052 13388
rect 6000 13345 6009 13379
rect 6009 13345 6043 13379
rect 6043 13345 6052 13379
rect 6000 13336 6052 13345
rect 9312 13336 9364 13388
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 10508 13379 10560 13388
rect 10508 13345 10517 13379
rect 10517 13345 10551 13379
rect 10551 13345 10560 13379
rect 10508 13336 10560 13345
rect 11520 13379 11572 13388
rect 11520 13345 11529 13379
rect 11529 13345 11563 13379
rect 11563 13345 11572 13379
rect 11520 13336 11572 13345
rect 10140 13268 10192 13320
rect 12348 13336 12400 13388
rect 11796 13268 11848 13320
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 14648 13336 14700 13388
rect 20076 13336 20128 13388
rect 13636 13268 13688 13320
rect 21732 13268 21784 13320
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 4620 13200 4672 13252
rect 4160 13132 4212 13184
rect 5908 13243 5960 13252
rect 5908 13209 5917 13243
rect 5917 13209 5951 13243
rect 5951 13209 5960 13243
rect 5908 13200 5960 13209
rect 10048 13200 10100 13252
rect 12072 13175 12124 13184
rect 12072 13141 12081 13175
rect 12081 13141 12115 13175
rect 12115 13141 12124 13175
rect 12072 13132 12124 13141
rect 13084 13200 13136 13252
rect 13360 13243 13412 13252
rect 13360 13209 13369 13243
rect 13369 13209 13403 13243
rect 13403 13209 13412 13243
rect 13360 13200 13412 13209
rect 12256 13132 12308 13184
rect 12808 13132 12860 13184
rect 19616 13132 19668 13184
rect 4266 13030 4318 13082
rect 4330 13030 4382 13082
rect 4394 13030 4446 13082
rect 4458 13030 4510 13082
rect 4522 13030 4574 13082
rect 9579 13030 9631 13082
rect 9643 13030 9695 13082
rect 9707 13030 9759 13082
rect 9771 13030 9823 13082
rect 9835 13030 9887 13082
rect 14892 13030 14944 13082
rect 14956 13030 15008 13082
rect 15020 13030 15072 13082
rect 15084 13030 15136 13082
rect 15148 13030 15200 13082
rect 20205 13030 20257 13082
rect 20269 13030 20321 13082
rect 20333 13030 20385 13082
rect 20397 13030 20449 13082
rect 20461 13030 20513 13082
rect 4160 12928 4212 12980
rect 4620 12928 4672 12980
rect 4712 12903 4764 12912
rect 4712 12869 4721 12903
rect 4721 12869 4755 12903
rect 4755 12869 4764 12903
rect 4712 12860 4764 12869
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 4896 12928 4948 12980
rect 12072 12928 12124 12980
rect 2872 12724 2924 12776
rect 4252 12724 4304 12776
rect 3148 12656 3200 12708
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5908 12792 5960 12844
rect 7196 12792 7248 12844
rect 12348 12860 12400 12912
rect 13084 12928 13136 12980
rect 21824 12928 21876 12980
rect 12256 12792 12308 12844
rect 12624 12835 12676 12844
rect 12624 12801 12633 12835
rect 12633 12801 12667 12835
rect 12667 12801 12676 12835
rect 13360 12860 13412 12912
rect 19340 12860 19392 12912
rect 19616 12903 19668 12912
rect 19616 12869 19625 12903
rect 19625 12869 19659 12903
rect 19659 12869 19668 12903
rect 19616 12860 19668 12869
rect 20536 12860 20588 12912
rect 12624 12792 12676 12801
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 5080 12699 5132 12708
rect 5080 12665 5089 12699
rect 5089 12665 5123 12699
rect 5123 12665 5132 12699
rect 5080 12656 5132 12665
rect 7656 12656 7708 12708
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 12808 12724 12860 12776
rect 18236 12767 18288 12776
rect 18236 12733 18245 12767
rect 18245 12733 18279 12767
rect 18279 12733 18288 12767
rect 18236 12724 18288 12733
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 15384 12656 15436 12708
rect 18052 12699 18104 12708
rect 18052 12665 18061 12699
rect 18061 12665 18095 12699
rect 18095 12665 18104 12699
rect 18052 12656 18104 12665
rect 18604 12656 18656 12708
rect 19432 12724 19484 12776
rect 19892 12767 19944 12776
rect 19892 12733 19901 12767
rect 19901 12733 19935 12767
rect 19935 12733 19944 12767
rect 19892 12724 19944 12733
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 15292 12588 15344 12640
rect 18420 12631 18472 12640
rect 18420 12597 18429 12631
rect 18429 12597 18463 12631
rect 18463 12597 18472 12631
rect 18420 12588 18472 12597
rect 18512 12631 18564 12640
rect 18512 12597 18521 12631
rect 18521 12597 18555 12631
rect 18555 12597 18564 12631
rect 18512 12588 18564 12597
rect 3606 12486 3658 12538
rect 3670 12486 3722 12538
rect 3734 12486 3786 12538
rect 3798 12486 3850 12538
rect 3862 12486 3914 12538
rect 8919 12486 8971 12538
rect 8983 12486 9035 12538
rect 9047 12486 9099 12538
rect 9111 12486 9163 12538
rect 9175 12486 9227 12538
rect 14232 12486 14284 12538
rect 14296 12486 14348 12538
rect 14360 12486 14412 12538
rect 14424 12486 14476 12538
rect 14488 12486 14540 12538
rect 19545 12486 19597 12538
rect 19609 12486 19661 12538
rect 19673 12486 19725 12538
rect 19737 12486 19789 12538
rect 19801 12486 19853 12538
rect 4252 12384 4304 12436
rect 4620 12384 4672 12436
rect 9404 12427 9456 12436
rect 9404 12393 9413 12427
rect 9413 12393 9447 12427
rect 9447 12393 9456 12427
rect 9404 12384 9456 12393
rect 12532 12384 12584 12436
rect 19432 12384 19484 12436
rect 20536 12384 20588 12436
rect 6920 12316 6972 12368
rect 14096 12316 14148 12368
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 8116 12248 8168 12300
rect 10416 12248 10468 12300
rect 17684 12248 17736 12300
rect 18236 12248 18288 12300
rect 18696 12291 18748 12300
rect 18696 12257 18705 12291
rect 18705 12257 18739 12291
rect 18739 12257 18748 12291
rect 18696 12248 18748 12257
rect 19892 12248 19944 12300
rect 4160 12180 4212 12232
rect 4712 12223 4764 12232
rect 4712 12189 4730 12223
rect 4730 12189 4764 12223
rect 4712 12180 4764 12189
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 12624 12223 12676 12232
rect 12624 12189 12658 12223
rect 12658 12189 12676 12223
rect 12624 12180 12676 12189
rect 8944 12112 8996 12164
rect 17040 12223 17092 12232
rect 17040 12189 17049 12223
rect 17049 12189 17083 12223
rect 17083 12189 17092 12223
rect 17040 12180 17092 12189
rect 18052 12180 18104 12232
rect 18512 12180 18564 12232
rect 19340 12180 19392 12232
rect 20444 12180 20496 12232
rect 17868 12112 17920 12164
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 7380 12087 7432 12096
rect 7380 12053 7389 12087
rect 7389 12053 7423 12087
rect 7423 12053 7432 12087
rect 7380 12044 7432 12053
rect 16948 12044 17000 12096
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 18328 12044 18380 12096
rect 4266 11942 4318 11994
rect 4330 11942 4382 11994
rect 4394 11942 4446 11994
rect 4458 11942 4510 11994
rect 4522 11942 4574 11994
rect 9579 11942 9631 11994
rect 9643 11942 9695 11994
rect 9707 11942 9759 11994
rect 9771 11942 9823 11994
rect 9835 11942 9887 11994
rect 14892 11942 14944 11994
rect 14956 11942 15008 11994
rect 15020 11942 15072 11994
rect 15084 11942 15136 11994
rect 15148 11942 15200 11994
rect 20205 11942 20257 11994
rect 20269 11942 20321 11994
rect 20333 11942 20385 11994
rect 20397 11942 20449 11994
rect 20461 11942 20513 11994
rect 6920 11840 6972 11892
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 17868 11840 17920 11892
rect 18328 11883 18380 11892
rect 18328 11849 18337 11883
rect 18337 11849 18371 11883
rect 18371 11849 18380 11883
rect 18328 11840 18380 11849
rect 848 11704 900 11756
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 1768 11704 1820 11756
rect 7012 11704 7064 11756
rect 7196 11636 7248 11688
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 10416 11704 10468 11756
rect 11336 11704 11388 11756
rect 10140 11636 10192 11688
rect 10968 11636 11020 11688
rect 7380 11568 7432 11620
rect 2228 11500 2280 11552
rect 6368 11500 6420 11552
rect 7104 11500 7156 11552
rect 8024 11568 8076 11620
rect 8576 11611 8628 11620
rect 8576 11577 8585 11611
rect 8585 11577 8619 11611
rect 8619 11577 8628 11611
rect 8576 11568 8628 11577
rect 10416 11568 10468 11620
rect 13820 11704 13872 11756
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 14004 11636 14056 11688
rect 18052 11772 18104 11824
rect 18236 11772 18288 11824
rect 18604 11772 18656 11824
rect 15844 11747 15896 11756
rect 15844 11713 15853 11747
rect 15853 11713 15887 11747
rect 15887 11713 15896 11747
rect 15844 11704 15896 11713
rect 15936 11704 15988 11756
rect 7656 11500 7708 11552
rect 9404 11500 9456 11552
rect 10600 11500 10652 11552
rect 12532 11500 12584 11552
rect 14556 11500 14608 11552
rect 14740 11500 14792 11552
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 16672 11543 16724 11552
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 16948 11636 17000 11688
rect 18144 11704 18196 11756
rect 22008 11747 22060 11756
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 18696 11636 18748 11688
rect 20628 11500 20680 11552
rect 3606 11398 3658 11450
rect 3670 11398 3722 11450
rect 3734 11398 3786 11450
rect 3798 11398 3850 11450
rect 3862 11398 3914 11450
rect 8919 11398 8971 11450
rect 8983 11398 9035 11450
rect 9047 11398 9099 11450
rect 9111 11398 9163 11450
rect 9175 11398 9227 11450
rect 14232 11398 14284 11450
rect 14296 11398 14348 11450
rect 14360 11398 14412 11450
rect 14424 11398 14476 11450
rect 14488 11398 14540 11450
rect 19545 11398 19597 11450
rect 19609 11398 19661 11450
rect 19673 11398 19725 11450
rect 19737 11398 19789 11450
rect 19801 11398 19853 11450
rect 8576 11296 8628 11348
rect 10416 11296 10468 11348
rect 15844 11296 15896 11348
rect 2688 11228 2740 11280
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 3332 11092 3384 11144
rect 5264 11160 5316 11212
rect 7012 11160 7064 11212
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 7288 11160 7340 11212
rect 10968 11228 11020 11280
rect 11336 11160 11388 11212
rect 11796 11203 11848 11212
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 12532 11203 12584 11212
rect 12532 11169 12541 11203
rect 12541 11169 12575 11203
rect 12575 11169 12584 11203
rect 12532 11160 12584 11169
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 7104 11092 7156 11144
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 13636 11160 13688 11212
rect 14004 11160 14056 11212
rect 14096 11160 14148 11212
rect 15384 11228 15436 11280
rect 16488 11228 16540 11280
rect 1952 11067 2004 11076
rect 1952 11033 1961 11067
rect 1961 11033 1995 11067
rect 1995 11033 2004 11067
rect 1952 11024 2004 11033
rect 3056 11067 3108 11076
rect 3056 11033 3065 11067
rect 3065 11033 3099 11067
rect 3099 11033 3108 11067
rect 3056 11024 3108 11033
rect 1768 10956 1820 11008
rect 2964 10956 3016 11008
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 3976 11024 4028 11076
rect 4712 11067 4764 11076
rect 4712 11033 4721 11067
rect 4721 11033 4755 11067
rect 4755 11033 4764 11067
rect 4712 11024 4764 11033
rect 6736 11024 6788 11076
rect 7840 11067 7892 11076
rect 7840 11033 7849 11067
rect 7849 11033 7883 11067
rect 7883 11033 7892 11067
rect 7840 11024 7892 11033
rect 8116 11024 8168 11076
rect 11796 11024 11848 11076
rect 12072 11024 12124 11076
rect 15936 11135 15988 11144
rect 15936 11101 15944 11135
rect 15944 11101 15988 11135
rect 15936 11092 15988 11101
rect 16212 11160 16264 11212
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 17684 11203 17736 11212
rect 17684 11169 17693 11203
rect 17693 11169 17727 11203
rect 17727 11169 17736 11203
rect 17684 11160 17736 11169
rect 4068 10956 4120 11008
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 10232 10999 10284 11008
rect 10232 10965 10241 10999
rect 10241 10965 10275 10999
rect 10275 10965 10284 10999
rect 10232 10956 10284 10965
rect 10692 10999 10744 11008
rect 10692 10965 10701 10999
rect 10701 10965 10735 10999
rect 10735 10965 10744 10999
rect 10692 10956 10744 10965
rect 11520 10999 11572 11008
rect 11520 10965 11529 10999
rect 11529 10965 11563 10999
rect 11563 10965 11572 10999
rect 11520 10956 11572 10965
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 11888 10956 11940 11008
rect 14464 10956 14516 11008
rect 15200 10956 15252 11008
rect 22008 11135 22060 11144
rect 22008 11101 22017 11135
rect 22017 11101 22051 11135
rect 22051 11101 22060 11135
rect 22008 11092 22060 11101
rect 18512 11024 18564 11076
rect 19064 10999 19116 11008
rect 19064 10965 19073 10999
rect 19073 10965 19107 10999
rect 19107 10965 19116 10999
rect 19064 10956 19116 10965
rect 4266 10854 4318 10906
rect 4330 10854 4382 10906
rect 4394 10854 4446 10906
rect 4458 10854 4510 10906
rect 4522 10854 4574 10906
rect 9579 10854 9631 10906
rect 9643 10854 9695 10906
rect 9707 10854 9759 10906
rect 9771 10854 9823 10906
rect 9835 10854 9887 10906
rect 14892 10854 14944 10906
rect 14956 10854 15008 10906
rect 15020 10854 15072 10906
rect 15084 10854 15136 10906
rect 15148 10854 15200 10906
rect 20205 10854 20257 10906
rect 20269 10854 20321 10906
rect 20333 10854 20385 10906
rect 20397 10854 20449 10906
rect 20461 10854 20513 10906
rect 2412 10727 2464 10736
rect 2412 10693 2421 10727
rect 2421 10693 2455 10727
rect 2455 10693 2464 10727
rect 2412 10684 2464 10693
rect 3240 10752 3292 10804
rect 5080 10752 5132 10804
rect 9036 10752 9088 10804
rect 11612 10752 11664 10804
rect 12072 10752 12124 10804
rect 16488 10752 16540 10804
rect 20720 10752 20772 10804
rect 3148 10616 3200 10668
rect 5816 10684 5868 10736
rect 3332 10616 3384 10668
rect 4528 10616 4580 10668
rect 2320 10591 2372 10600
rect 2320 10557 2329 10591
rect 2329 10557 2363 10591
rect 2363 10557 2372 10591
rect 2320 10548 2372 10557
rect 2964 10591 3016 10600
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 3424 10548 3476 10600
rect 4068 10548 4120 10600
rect 7380 10684 7432 10736
rect 7840 10684 7892 10736
rect 10232 10684 10284 10736
rect 11336 10727 11388 10736
rect 11336 10693 11345 10727
rect 11345 10693 11379 10727
rect 11379 10693 11388 10727
rect 11336 10684 11388 10693
rect 6736 10616 6788 10668
rect 3056 10480 3108 10532
rect 4988 10480 5040 10532
rect 7196 10616 7248 10668
rect 11612 10616 11664 10668
rect 11888 10659 11940 10668
rect 11888 10625 11932 10659
rect 11932 10625 11940 10659
rect 11888 10616 11940 10625
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 15292 10684 15344 10736
rect 14740 10616 14792 10668
rect 14004 10548 14056 10557
rect 14556 10591 14608 10600
rect 14556 10557 14565 10591
rect 14565 10557 14599 10591
rect 14599 10557 14608 10591
rect 14556 10548 14608 10557
rect 19340 10616 19392 10668
rect 20444 10616 20496 10668
rect 7564 10480 7616 10532
rect 3332 10412 3384 10464
rect 4160 10412 4212 10464
rect 4896 10412 4948 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 8208 10412 8260 10464
rect 13820 10523 13872 10532
rect 13820 10489 13829 10523
rect 13829 10489 13863 10523
rect 13863 10489 13872 10523
rect 13820 10480 13872 10489
rect 14464 10480 14516 10532
rect 15476 10480 15528 10532
rect 19984 10480 20036 10532
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 11980 10412 12032 10464
rect 14096 10412 14148 10464
rect 14648 10412 14700 10464
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 19432 10412 19484 10464
rect 20076 10455 20128 10464
rect 20076 10421 20085 10455
rect 20085 10421 20119 10455
rect 20119 10421 20128 10455
rect 20076 10412 20128 10421
rect 20536 10412 20588 10464
rect 3606 10310 3658 10362
rect 3670 10310 3722 10362
rect 3734 10310 3786 10362
rect 3798 10310 3850 10362
rect 3862 10310 3914 10362
rect 8919 10310 8971 10362
rect 8983 10310 9035 10362
rect 9047 10310 9099 10362
rect 9111 10310 9163 10362
rect 9175 10310 9227 10362
rect 14232 10310 14284 10362
rect 14296 10310 14348 10362
rect 14360 10310 14412 10362
rect 14424 10310 14476 10362
rect 14488 10310 14540 10362
rect 19545 10310 19597 10362
rect 19609 10310 19661 10362
rect 19673 10310 19725 10362
rect 19737 10310 19789 10362
rect 19801 10310 19853 10362
rect 2320 10208 2372 10260
rect 3976 10208 4028 10260
rect 4528 10251 4580 10260
rect 4528 10217 4537 10251
rect 4537 10217 4571 10251
rect 4571 10217 4580 10251
rect 4528 10208 4580 10217
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 2228 10115 2280 10124
rect 2228 10081 2237 10115
rect 2237 10081 2271 10115
rect 2271 10081 2280 10115
rect 2228 10072 2280 10081
rect 3332 10140 3384 10192
rect 4160 10140 4212 10192
rect 5816 10208 5868 10260
rect 8116 10208 8168 10260
rect 10692 10208 10744 10260
rect 13176 10208 13228 10260
rect 15384 10208 15436 10260
rect 18696 10208 18748 10260
rect 19524 10208 19576 10260
rect 19984 10208 20036 10260
rect 3424 10072 3476 10124
rect 4896 10115 4948 10124
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 4896 10072 4948 10081
rect 1768 10004 1820 10056
rect 2412 10004 2464 10056
rect 4620 10004 4672 10056
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 7196 10072 7248 10124
rect 6736 10004 6788 10056
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10968 10004 11020 10056
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 6276 9936 6328 9988
rect 12348 10047 12400 10056
rect 12348 10013 12357 10047
rect 12357 10013 12391 10047
rect 12391 10013 12400 10047
rect 12348 10004 12400 10013
rect 15568 10140 15620 10192
rect 21180 10140 21232 10192
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 12900 10004 12952 10056
rect 6460 9911 6512 9920
rect 6460 9877 6469 9911
rect 6469 9877 6503 9911
rect 6503 9877 6512 9911
rect 6460 9868 6512 9877
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 13268 9936 13320 9988
rect 15292 10072 15344 10124
rect 16948 10072 17000 10124
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 16672 10004 16724 10056
rect 17868 10004 17920 10056
rect 18420 10072 18472 10124
rect 19064 10072 19116 10124
rect 19432 10072 19484 10124
rect 18696 10004 18748 10056
rect 20536 10115 20588 10124
rect 20536 10081 20545 10115
rect 20545 10081 20579 10115
rect 20579 10081 20588 10115
rect 20536 10072 20588 10081
rect 20628 10115 20680 10124
rect 20628 10081 20637 10115
rect 20637 10081 20671 10115
rect 20671 10081 20680 10115
rect 20628 10072 20680 10081
rect 20720 10072 20772 10124
rect 20444 10047 20496 10056
rect 20444 10013 20453 10047
rect 20453 10013 20487 10047
rect 20487 10013 20496 10047
rect 20444 10004 20496 10013
rect 21732 10047 21784 10056
rect 21732 10013 21741 10047
rect 21741 10013 21775 10047
rect 21775 10013 21784 10047
rect 21732 10004 21784 10013
rect 15384 9936 15436 9988
rect 14556 9868 14608 9920
rect 14648 9868 14700 9920
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 18052 9911 18104 9920
rect 18052 9877 18061 9911
rect 18061 9877 18095 9911
rect 18095 9877 18104 9911
rect 18052 9868 18104 9877
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 18880 9868 18932 9920
rect 19616 9911 19668 9920
rect 19616 9877 19625 9911
rect 19625 9877 19659 9911
rect 19659 9877 19668 9911
rect 19616 9868 19668 9877
rect 20628 9868 20680 9920
rect 21272 9911 21324 9920
rect 21272 9877 21281 9911
rect 21281 9877 21315 9911
rect 21315 9877 21324 9911
rect 21272 9868 21324 9877
rect 21364 9911 21416 9920
rect 21364 9877 21373 9911
rect 21373 9877 21407 9911
rect 21407 9877 21416 9911
rect 21364 9868 21416 9877
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 4266 9766 4318 9818
rect 4330 9766 4382 9818
rect 4394 9766 4446 9818
rect 4458 9766 4510 9818
rect 4522 9766 4574 9818
rect 9579 9766 9631 9818
rect 9643 9766 9695 9818
rect 9707 9766 9759 9818
rect 9771 9766 9823 9818
rect 9835 9766 9887 9818
rect 14892 9766 14944 9818
rect 14956 9766 15008 9818
rect 15020 9766 15072 9818
rect 15084 9766 15136 9818
rect 15148 9766 15200 9818
rect 20205 9766 20257 9818
rect 20269 9766 20321 9818
rect 20333 9766 20385 9818
rect 20397 9766 20449 9818
rect 20461 9766 20513 9818
rect 2136 9664 2188 9716
rect 7564 9664 7616 9716
rect 12716 9664 12768 9716
rect 19616 9664 19668 9716
rect 21364 9664 21416 9716
rect 4712 9596 4764 9648
rect 12808 9596 12860 9648
rect 15384 9596 15436 9648
rect 4160 9528 4212 9580
rect 6736 9528 6788 9580
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 14740 9528 14792 9580
rect 16856 9596 16908 9648
rect 16764 9571 16816 9580
rect 16764 9537 16773 9571
rect 16773 9537 16807 9571
rect 16807 9537 16816 9571
rect 16764 9528 16816 9537
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 17868 9571 17920 9580
rect 17868 9537 17877 9571
rect 17877 9537 17911 9571
rect 17911 9537 17920 9571
rect 17868 9528 17920 9537
rect 18144 9528 18196 9580
rect 18880 9571 18932 9580
rect 18880 9537 18889 9571
rect 18889 9537 18923 9571
rect 18923 9537 18932 9571
rect 18880 9528 18932 9537
rect 4620 9460 4672 9512
rect 18052 9460 18104 9512
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 4160 9392 4212 9444
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 19892 9528 19944 9580
rect 20168 9639 20220 9648
rect 20168 9605 20177 9639
rect 20177 9605 20211 9639
rect 20211 9605 20220 9639
rect 20168 9596 20220 9605
rect 21732 9596 21784 9648
rect 21272 9528 21324 9580
rect 19340 9460 19392 9512
rect 20628 9460 20680 9512
rect 15568 9324 15620 9376
rect 19984 9324 20036 9376
rect 3606 9222 3658 9274
rect 3670 9222 3722 9274
rect 3734 9222 3786 9274
rect 3798 9222 3850 9274
rect 3862 9222 3914 9274
rect 8919 9222 8971 9274
rect 8983 9222 9035 9274
rect 9047 9222 9099 9274
rect 9111 9222 9163 9274
rect 9175 9222 9227 9274
rect 14232 9222 14284 9274
rect 14296 9222 14348 9274
rect 14360 9222 14412 9274
rect 14424 9222 14476 9274
rect 14488 9222 14540 9274
rect 19545 9222 19597 9274
rect 19609 9222 19661 9274
rect 19673 9222 19725 9274
rect 19737 9222 19789 9274
rect 19801 9222 19853 9274
rect 848 9052 900 9104
rect 6460 9120 6512 9172
rect 6736 9163 6788 9172
rect 6736 9129 6745 9163
rect 6745 9129 6779 9163
rect 6779 9129 6788 9163
rect 6736 9120 6788 9129
rect 19892 9120 19944 9172
rect 1676 8780 1728 8832
rect 9404 9052 9456 9104
rect 5816 8984 5868 9036
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 7380 9027 7432 9036
rect 7380 8993 7389 9027
rect 7389 8993 7423 9027
rect 7423 8993 7432 9027
rect 7380 8984 7432 8993
rect 7288 8916 7340 8968
rect 7748 8916 7800 8968
rect 11520 8984 11572 9036
rect 15292 9052 15344 9104
rect 15384 9052 15436 9104
rect 9496 8848 9548 8900
rect 10324 8959 10376 8968
rect 10324 8925 10368 8959
rect 10368 8925 10376 8959
rect 10324 8916 10376 8925
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 12532 8959 12584 8968
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 12716 8916 12768 8968
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 18420 9095 18472 9104
rect 18420 9061 18429 9095
rect 18429 9061 18463 9095
rect 18463 9061 18472 9095
rect 18420 9052 18472 9061
rect 15476 8959 15528 8968
rect 15476 8925 15485 8959
rect 15485 8925 15519 8959
rect 15519 8925 15528 8959
rect 15476 8916 15528 8925
rect 16764 8984 16816 9036
rect 18788 8984 18840 9036
rect 6920 8780 6972 8832
rect 10416 8780 10468 8832
rect 21916 8823 21968 8832
rect 21916 8789 21925 8823
rect 21925 8789 21959 8823
rect 21959 8789 21968 8823
rect 21916 8780 21968 8789
rect 4266 8678 4318 8730
rect 4330 8678 4382 8730
rect 4394 8678 4446 8730
rect 4458 8678 4510 8730
rect 4522 8678 4574 8730
rect 9579 8678 9631 8730
rect 9643 8678 9695 8730
rect 9707 8678 9759 8730
rect 9771 8678 9823 8730
rect 9835 8678 9887 8730
rect 14892 8678 14944 8730
rect 14956 8678 15008 8730
rect 15020 8678 15072 8730
rect 15084 8678 15136 8730
rect 15148 8678 15200 8730
rect 20205 8678 20257 8730
rect 20269 8678 20321 8730
rect 20333 8678 20385 8730
rect 20397 8678 20449 8730
rect 20461 8678 20513 8730
rect 4160 8576 4212 8628
rect 9496 8576 9548 8628
rect 4344 8508 4396 8560
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 3056 8440 3108 8492
rect 4068 8483 4120 8492
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 4160 8440 4212 8492
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 10232 8508 10284 8560
rect 9588 8440 9640 8492
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 3240 8347 3292 8356
rect 3240 8313 3249 8347
rect 3249 8313 3283 8347
rect 3283 8313 3292 8347
rect 3240 8304 3292 8313
rect 4252 8304 4304 8356
rect 5540 8304 5592 8356
rect 7104 8304 7156 8356
rect 5632 8279 5684 8288
rect 5632 8245 5641 8279
rect 5641 8245 5675 8279
rect 5675 8245 5684 8279
rect 5632 8236 5684 8245
rect 9312 8372 9364 8424
rect 9404 8372 9456 8424
rect 10600 8440 10652 8492
rect 11520 8551 11572 8560
rect 11520 8517 11529 8551
rect 11529 8517 11563 8551
rect 11563 8517 11572 8551
rect 11520 8508 11572 8517
rect 12716 8551 12768 8560
rect 12716 8517 12725 8551
rect 12725 8517 12759 8551
rect 12759 8517 12768 8551
rect 12716 8508 12768 8517
rect 12624 8440 12676 8492
rect 13268 8440 13320 8492
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 15292 8440 15344 8492
rect 17132 8440 17184 8492
rect 19984 8483 20036 8492
rect 11244 8372 11296 8424
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 19248 8372 19300 8424
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 9588 8304 9640 8356
rect 16212 8304 16264 8356
rect 21548 8347 21600 8356
rect 21548 8313 21557 8347
rect 21557 8313 21591 8347
rect 21591 8313 21600 8347
rect 21548 8304 21600 8313
rect 9404 8236 9456 8288
rect 17592 8279 17644 8288
rect 17592 8245 17601 8279
rect 17601 8245 17635 8279
rect 17635 8245 17644 8279
rect 17592 8236 17644 8245
rect 18972 8279 19024 8288
rect 18972 8245 18981 8279
rect 18981 8245 19015 8279
rect 19015 8245 19024 8279
rect 18972 8236 19024 8245
rect 19432 8236 19484 8288
rect 3606 8134 3658 8186
rect 3670 8134 3722 8186
rect 3734 8134 3786 8186
rect 3798 8134 3850 8186
rect 3862 8134 3914 8186
rect 8919 8134 8971 8186
rect 8983 8134 9035 8186
rect 9047 8134 9099 8186
rect 9111 8134 9163 8186
rect 9175 8134 9227 8186
rect 14232 8134 14284 8186
rect 14296 8134 14348 8186
rect 14360 8134 14412 8186
rect 14424 8134 14476 8186
rect 14488 8134 14540 8186
rect 19545 8134 19597 8186
rect 19609 8134 19661 8186
rect 19673 8134 19725 8186
rect 19737 8134 19789 8186
rect 19801 8134 19853 8186
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 4068 8032 4120 8084
rect 9312 8032 9364 8084
rect 12256 8032 12308 8084
rect 12532 8032 12584 8084
rect 1952 7896 2004 7948
rect 3240 7896 3292 7948
rect 5448 7964 5500 8016
rect 4344 7896 4396 7948
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 12440 7964 12492 8016
rect 9588 7939 9640 7948
rect 4252 7828 4304 7880
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 6828 7828 6880 7880
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 7656 7828 7708 7880
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 9404 7828 9456 7880
rect 9588 7905 9597 7939
rect 9597 7905 9631 7939
rect 9631 7905 9640 7939
rect 9588 7896 9640 7905
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 13268 7896 13320 7905
rect 14004 7896 14056 7948
rect 14556 7939 14608 7948
rect 14556 7905 14565 7939
rect 14565 7905 14599 7939
rect 14599 7905 14608 7939
rect 14556 7896 14608 7905
rect 16948 7939 17000 7948
rect 16948 7905 16957 7939
rect 16957 7905 16991 7939
rect 16991 7905 17000 7939
rect 16948 7896 17000 7905
rect 17592 7896 17644 7948
rect 4620 7760 4672 7812
rect 8392 7760 8444 7812
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 10600 7871 10652 7880
rect 10600 7837 10609 7871
rect 10609 7837 10643 7871
rect 10643 7837 10652 7871
rect 10600 7828 10652 7837
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 14832 7871 14884 7880
rect 14832 7837 14841 7871
rect 14841 7837 14875 7871
rect 14875 7837 14884 7871
rect 14832 7828 14884 7837
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 1768 7735 1820 7744
rect 1768 7701 1777 7735
rect 1777 7701 1811 7735
rect 1811 7701 1820 7735
rect 1768 7692 1820 7701
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 2596 7735 2648 7744
rect 2596 7701 2605 7735
rect 2605 7701 2639 7735
rect 2639 7701 2648 7735
rect 2596 7692 2648 7701
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 5080 7692 5132 7744
rect 5356 7692 5408 7744
rect 5540 7692 5592 7744
rect 7380 7735 7432 7744
rect 7380 7701 7389 7735
rect 7389 7701 7423 7735
rect 7423 7701 7432 7735
rect 7380 7692 7432 7701
rect 9956 7735 10008 7744
rect 9956 7701 9965 7735
rect 9965 7701 9999 7735
rect 9999 7701 10008 7735
rect 9956 7692 10008 7701
rect 10140 7692 10192 7744
rect 12992 7735 13044 7744
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 13084 7735 13136 7744
rect 13084 7701 13093 7735
rect 13093 7701 13127 7735
rect 13127 7701 13136 7735
rect 13084 7692 13136 7701
rect 15292 7692 15344 7744
rect 17224 7828 17276 7880
rect 17868 7828 17920 7880
rect 19248 7896 19300 7948
rect 19432 7828 19484 7880
rect 18144 7760 18196 7812
rect 19616 7735 19668 7744
rect 19616 7701 19625 7735
rect 19625 7701 19659 7735
rect 19659 7701 19668 7735
rect 19616 7692 19668 7701
rect 19892 7692 19944 7744
rect 21916 7735 21968 7744
rect 21916 7701 21925 7735
rect 21925 7701 21959 7735
rect 21959 7701 21968 7735
rect 21916 7692 21968 7701
rect 4266 7590 4318 7642
rect 4330 7590 4382 7642
rect 4394 7590 4446 7642
rect 4458 7590 4510 7642
rect 4522 7590 4574 7642
rect 9579 7590 9631 7642
rect 9643 7590 9695 7642
rect 9707 7590 9759 7642
rect 9771 7590 9823 7642
rect 9835 7590 9887 7642
rect 14892 7590 14944 7642
rect 14956 7590 15008 7642
rect 15020 7590 15072 7642
rect 15084 7590 15136 7642
rect 15148 7590 15200 7642
rect 20205 7590 20257 7642
rect 20269 7590 20321 7642
rect 20333 7590 20385 7642
rect 20397 7590 20449 7642
rect 20461 7590 20513 7642
rect 1768 7488 1820 7540
rect 2596 7488 2648 7540
rect 5356 7531 5408 7540
rect 5356 7497 5365 7531
rect 5365 7497 5399 7531
rect 5399 7497 5408 7531
rect 5356 7488 5408 7497
rect 7196 7488 7248 7540
rect 12992 7488 13044 7540
rect 19616 7488 19668 7540
rect 2412 7420 2464 7472
rect 4160 7420 4212 7472
rect 5080 7420 5132 7472
rect 9956 7463 10008 7472
rect 9956 7429 9965 7463
rect 9965 7429 9999 7463
rect 9999 7429 10008 7463
rect 9956 7420 10008 7429
rect 10140 7463 10192 7472
rect 10140 7429 10149 7463
rect 10149 7429 10183 7463
rect 10183 7429 10192 7463
rect 10140 7420 10192 7429
rect 13084 7420 13136 7472
rect 18972 7420 19024 7472
rect 848 7352 900 7404
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 1860 7352 1912 7404
rect 2596 7395 2648 7404
rect 2596 7361 2640 7395
rect 2640 7361 2648 7395
rect 2596 7352 2648 7361
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 3056 7284 3108 7336
rect 4712 7352 4764 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 4804 7284 4856 7336
rect 6000 7284 6052 7336
rect 12532 7395 12584 7404
rect 12532 7361 12541 7395
rect 12541 7361 12575 7395
rect 12575 7361 12584 7395
rect 12532 7352 12584 7361
rect 14096 7352 14148 7404
rect 14740 7352 14792 7404
rect 15200 7352 15252 7404
rect 19340 7420 19392 7472
rect 1860 7259 1912 7268
rect 1860 7225 1869 7259
rect 1869 7225 1903 7259
rect 1903 7225 1912 7259
rect 1860 7216 1912 7225
rect 1952 7216 2004 7268
rect 4160 7216 4212 7268
rect 12348 7216 12400 7268
rect 16764 7216 16816 7268
rect 19248 7327 19300 7336
rect 19248 7293 19257 7327
rect 19257 7293 19291 7327
rect 19291 7293 19300 7327
rect 19248 7284 19300 7293
rect 19432 7216 19484 7268
rect 19984 7284 20036 7336
rect 20536 7284 20588 7336
rect 21824 7352 21876 7404
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 20260 7259 20312 7268
rect 20260 7225 20269 7259
rect 20269 7225 20303 7259
rect 20303 7225 20312 7259
rect 20260 7216 20312 7225
rect 7840 7191 7892 7200
rect 7840 7157 7849 7191
rect 7849 7157 7883 7191
rect 7883 7157 7892 7191
rect 7840 7148 7892 7157
rect 10324 7191 10376 7200
rect 10324 7157 10333 7191
rect 10333 7157 10367 7191
rect 10367 7157 10376 7191
rect 10324 7148 10376 7157
rect 15568 7148 15620 7200
rect 18328 7191 18380 7200
rect 18328 7157 18337 7191
rect 18337 7157 18371 7191
rect 18371 7157 18380 7191
rect 18328 7148 18380 7157
rect 20904 7148 20956 7200
rect 3606 7046 3658 7098
rect 3670 7046 3722 7098
rect 3734 7046 3786 7098
rect 3798 7046 3850 7098
rect 3862 7046 3914 7098
rect 8919 7046 8971 7098
rect 8983 7046 9035 7098
rect 9047 7046 9099 7098
rect 9111 7046 9163 7098
rect 9175 7046 9227 7098
rect 14232 7046 14284 7098
rect 14296 7046 14348 7098
rect 14360 7046 14412 7098
rect 14424 7046 14476 7098
rect 14488 7046 14540 7098
rect 19545 7046 19597 7098
rect 19609 7046 19661 7098
rect 19673 7046 19725 7098
rect 19737 7046 19789 7098
rect 19801 7046 19853 7098
rect 6828 6944 6880 6996
rect 15200 6944 15252 6996
rect 19892 6987 19944 6996
rect 19892 6953 19901 6987
rect 19901 6953 19935 6987
rect 19935 6953 19944 6987
rect 19892 6944 19944 6953
rect 17224 6876 17276 6928
rect 5264 6808 5316 6860
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 6552 6808 6604 6860
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 14648 6808 14700 6860
rect 15844 6808 15896 6860
rect 16120 6851 16172 6860
rect 16120 6817 16129 6851
rect 16129 6817 16163 6851
rect 16163 6817 16172 6851
rect 16120 6808 16172 6817
rect 16948 6808 17000 6860
rect 18328 6808 18380 6860
rect 19064 6808 19116 6860
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 5080 6715 5132 6724
rect 5080 6681 5089 6715
rect 5089 6681 5123 6715
rect 5123 6681 5132 6715
rect 5080 6672 5132 6681
rect 5264 6672 5316 6724
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 13912 6740 13964 6792
rect 20720 6876 20772 6928
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 19432 6740 19484 6792
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 20260 6783 20312 6792
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 20536 6740 20588 6792
rect 16580 6672 16632 6724
rect 18236 6672 18288 6724
rect 3332 6604 3384 6656
rect 5540 6604 5592 6656
rect 6092 6647 6144 6656
rect 6092 6613 6101 6647
rect 6101 6613 6135 6647
rect 6135 6613 6144 6647
rect 6092 6604 6144 6613
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 16672 6604 16724 6656
rect 17132 6604 17184 6656
rect 18420 6604 18472 6656
rect 18788 6604 18840 6656
rect 21824 6604 21876 6656
rect 4266 6502 4318 6554
rect 4330 6502 4382 6554
rect 4394 6502 4446 6554
rect 4458 6502 4510 6554
rect 4522 6502 4574 6554
rect 9579 6502 9631 6554
rect 9643 6502 9695 6554
rect 9707 6502 9759 6554
rect 9771 6502 9823 6554
rect 9835 6502 9887 6554
rect 14892 6502 14944 6554
rect 14956 6502 15008 6554
rect 15020 6502 15072 6554
rect 15084 6502 15136 6554
rect 15148 6502 15200 6554
rect 20205 6502 20257 6554
rect 20269 6502 20321 6554
rect 20333 6502 20385 6554
rect 20397 6502 20449 6554
rect 20461 6502 20513 6554
rect 2596 6400 2648 6452
rect 4804 6400 4856 6452
rect 5264 6443 5316 6452
rect 5264 6409 5273 6443
rect 5273 6409 5307 6443
rect 5307 6409 5316 6443
rect 5264 6400 5316 6409
rect 6092 6400 6144 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 7656 6400 7708 6452
rect 8392 6400 8444 6452
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 19340 6400 19392 6452
rect 4988 6332 5040 6384
rect 5448 6375 5500 6384
rect 5448 6341 5457 6375
rect 5457 6341 5491 6375
rect 5491 6341 5500 6375
rect 5448 6332 5500 6341
rect 14648 6375 14700 6384
rect 14648 6341 14657 6375
rect 14657 6341 14691 6375
rect 14691 6341 14700 6375
rect 14648 6332 14700 6341
rect 16120 6332 16172 6384
rect 848 6264 900 6316
rect 3516 6264 3568 6316
rect 3976 6264 4028 6316
rect 4160 6264 4212 6316
rect 6092 6264 6144 6316
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 9496 6264 9548 6316
rect 9772 6264 9824 6316
rect 12072 6264 12124 6316
rect 12348 6307 12400 6316
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 4712 6239 4764 6248
rect 4712 6205 4721 6239
rect 4721 6205 4755 6239
rect 4755 6205 4764 6239
rect 4712 6196 4764 6205
rect 5356 6196 5408 6248
rect 7012 6239 7064 6248
rect 7012 6205 7021 6239
rect 7021 6205 7055 6239
rect 7055 6205 7064 6239
rect 7012 6196 7064 6205
rect 4896 6128 4948 6180
rect 6552 6128 6604 6180
rect 7564 6239 7616 6248
rect 7564 6205 7573 6239
rect 7573 6205 7607 6239
rect 7607 6205 7616 6239
rect 7564 6196 7616 6205
rect 9404 6239 9456 6248
rect 9404 6205 9413 6239
rect 9413 6205 9447 6239
rect 9447 6205 9456 6239
rect 9404 6196 9456 6205
rect 10232 6239 10284 6248
rect 10232 6205 10241 6239
rect 10241 6205 10275 6239
rect 10275 6205 10284 6239
rect 10232 6196 10284 6205
rect 13084 6264 13136 6316
rect 13820 6264 13872 6316
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 20076 6307 20128 6316
rect 20076 6273 20085 6307
rect 20085 6273 20119 6307
rect 20119 6273 20128 6307
rect 20076 6264 20128 6273
rect 21180 6264 21232 6316
rect 12072 6171 12124 6180
rect 12072 6137 12081 6171
rect 12081 6137 12115 6171
rect 12115 6137 12124 6171
rect 12072 6128 12124 6137
rect 13912 6196 13964 6248
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 18880 6239 18932 6248
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 20536 6196 20588 6248
rect 12532 6128 12584 6180
rect 14096 6128 14148 6180
rect 4068 6060 4120 6112
rect 4804 6060 4856 6112
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 12992 6060 13044 6112
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 18788 6128 18840 6180
rect 21548 6171 21600 6180
rect 21548 6137 21557 6171
rect 21557 6137 21591 6171
rect 21591 6137 21600 6171
rect 21548 6128 21600 6137
rect 14924 6103 14976 6112
rect 14924 6069 14933 6103
rect 14933 6069 14967 6103
rect 14967 6069 14976 6103
rect 14924 6060 14976 6069
rect 3606 5958 3658 6010
rect 3670 5958 3722 6010
rect 3734 5958 3786 6010
rect 3798 5958 3850 6010
rect 3862 5958 3914 6010
rect 8919 5958 8971 6010
rect 8983 5958 9035 6010
rect 9047 5958 9099 6010
rect 9111 5958 9163 6010
rect 9175 5958 9227 6010
rect 14232 5958 14284 6010
rect 14296 5958 14348 6010
rect 14360 5958 14412 6010
rect 14424 5958 14476 6010
rect 14488 5958 14540 6010
rect 19545 5958 19597 6010
rect 19609 5958 19661 6010
rect 19673 5958 19725 6010
rect 19737 5958 19789 6010
rect 19801 5958 19853 6010
rect 3976 5856 4028 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 7564 5899 7616 5908
rect 7564 5865 7573 5899
rect 7573 5865 7607 5899
rect 7607 5865 7616 5899
rect 7564 5856 7616 5865
rect 8116 5856 8168 5908
rect 9772 5899 9824 5908
rect 9772 5865 9781 5899
rect 9781 5865 9815 5899
rect 9815 5865 9824 5899
rect 9772 5856 9824 5865
rect 10692 5899 10744 5908
rect 10692 5865 10701 5899
rect 10701 5865 10735 5899
rect 10735 5865 10744 5899
rect 10692 5856 10744 5865
rect 12532 5856 12584 5908
rect 14648 5856 14700 5908
rect 21824 5899 21876 5908
rect 21824 5865 21833 5899
rect 21833 5865 21867 5899
rect 21867 5865 21876 5899
rect 21824 5856 21876 5865
rect 4252 5720 4304 5772
rect 3332 5652 3384 5704
rect 3976 5652 4028 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 4620 5652 4672 5704
rect 5448 5720 5500 5772
rect 10232 5788 10284 5840
rect 14004 5788 14056 5840
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 7012 5652 7064 5704
rect 7196 5652 7248 5704
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 10324 5720 10376 5772
rect 11796 5720 11848 5772
rect 14924 5763 14976 5772
rect 14924 5729 14933 5763
rect 14933 5729 14967 5763
rect 14967 5729 14976 5763
rect 14924 5720 14976 5729
rect 19064 5831 19116 5840
rect 19064 5797 19073 5831
rect 19073 5797 19107 5831
rect 19107 5797 19116 5831
rect 19064 5788 19116 5797
rect 10048 5584 10100 5636
rect 12072 5652 12124 5704
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 13176 5695 13228 5704
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 22008 5695 22060 5704
rect 22008 5661 22017 5695
rect 22017 5661 22051 5695
rect 22051 5661 22060 5695
rect 22008 5652 22060 5661
rect 12532 5584 12584 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 4068 5516 4120 5568
rect 4252 5516 4304 5568
rect 7564 5516 7616 5568
rect 7932 5559 7984 5568
rect 7932 5525 7941 5559
rect 7941 5525 7975 5559
rect 7975 5525 7984 5559
rect 7932 5516 7984 5525
rect 11796 5516 11848 5568
rect 13820 5516 13872 5568
rect 14740 5516 14792 5568
rect 18696 5559 18748 5568
rect 18696 5525 18705 5559
rect 18705 5525 18739 5559
rect 18739 5525 18748 5559
rect 18696 5516 18748 5525
rect 4266 5414 4318 5466
rect 4330 5414 4382 5466
rect 4394 5414 4446 5466
rect 4458 5414 4510 5466
rect 4522 5414 4574 5466
rect 9579 5414 9631 5466
rect 9643 5414 9695 5466
rect 9707 5414 9759 5466
rect 9771 5414 9823 5466
rect 9835 5414 9887 5466
rect 14892 5414 14944 5466
rect 14956 5414 15008 5466
rect 15020 5414 15072 5466
rect 15084 5414 15136 5466
rect 15148 5414 15200 5466
rect 20205 5414 20257 5466
rect 20269 5414 20321 5466
rect 20333 5414 20385 5466
rect 20397 5414 20449 5466
rect 20461 5414 20513 5466
rect 3516 5312 3568 5364
rect 4068 5312 4120 5364
rect 4160 5312 4212 5364
rect 4804 5312 4856 5364
rect 11796 5312 11848 5364
rect 12348 5312 12400 5364
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 21272 5312 21324 5364
rect 848 5176 900 5228
rect 4620 5244 4672 5296
rect 4988 5287 5040 5296
rect 4988 5253 4997 5287
rect 4997 5253 5031 5287
rect 5031 5253 5040 5287
rect 4988 5244 5040 5253
rect 10692 5244 10744 5296
rect 17224 5244 17276 5296
rect 3976 5108 4028 5160
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 5724 5108 5776 5160
rect 7288 5108 7340 5160
rect 7932 5151 7984 5160
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 14096 5176 14148 5228
rect 15108 5176 15160 5228
rect 11980 5108 12032 5160
rect 13728 5108 13780 5160
rect 14648 5108 14700 5160
rect 16672 5108 16724 5160
rect 17040 5108 17092 5160
rect 17684 5176 17736 5228
rect 17868 5151 17920 5160
rect 17868 5117 17877 5151
rect 17877 5117 17911 5151
rect 17911 5117 17920 5151
rect 17868 5108 17920 5117
rect 19156 5176 19208 5228
rect 22008 5219 22060 5228
rect 22008 5185 22017 5219
rect 22017 5185 22051 5219
rect 22051 5185 22060 5219
rect 22008 5176 22060 5185
rect 18880 5108 18932 5160
rect 19340 5151 19392 5160
rect 19340 5117 19349 5151
rect 19349 5117 19383 5151
rect 19383 5117 19392 5151
rect 19340 5108 19392 5117
rect 19248 5040 19300 5092
rect 3606 4870 3658 4922
rect 3670 4870 3722 4922
rect 3734 4870 3786 4922
rect 3798 4870 3850 4922
rect 3862 4870 3914 4922
rect 8919 4870 8971 4922
rect 8983 4870 9035 4922
rect 9047 4870 9099 4922
rect 9111 4870 9163 4922
rect 9175 4870 9227 4922
rect 14232 4870 14284 4922
rect 14296 4870 14348 4922
rect 14360 4870 14412 4922
rect 14424 4870 14476 4922
rect 14488 4870 14540 4922
rect 19545 4870 19597 4922
rect 19609 4870 19661 4922
rect 19673 4870 19725 4922
rect 19737 4870 19789 4922
rect 19801 4870 19853 4922
rect 5080 4768 5132 4820
rect 9588 4768 9640 4820
rect 10048 4768 10100 4820
rect 13912 4811 13964 4820
rect 13912 4777 13921 4811
rect 13921 4777 13955 4811
rect 13955 4777 13964 4811
rect 13912 4768 13964 4777
rect 14740 4768 14792 4820
rect 17684 4811 17736 4820
rect 17684 4777 17693 4811
rect 17693 4777 17727 4811
rect 17727 4777 17736 4811
rect 17684 4768 17736 4777
rect 17868 4768 17920 4820
rect 19248 4811 19300 4820
rect 19248 4777 19257 4811
rect 19257 4777 19291 4811
rect 19291 4777 19300 4811
rect 19248 4768 19300 4777
rect 9496 4743 9548 4752
rect 9496 4709 9505 4743
rect 9505 4709 9539 4743
rect 9539 4709 9548 4743
rect 9496 4700 9548 4709
rect 4712 4632 4764 4684
rect 848 4564 900 4616
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 9404 4675 9456 4684
rect 9404 4641 9413 4675
rect 9413 4641 9447 4675
rect 9447 4641 9456 4675
rect 9404 4632 9456 4641
rect 10232 4632 10284 4684
rect 10784 4675 10836 4684
rect 6920 4564 6972 4616
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 14648 4632 14700 4684
rect 19156 4700 19208 4752
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 7748 4496 7800 4548
rect 10140 4496 10192 4548
rect 13544 4539 13596 4548
rect 13544 4505 13553 4539
rect 13553 4505 13587 4539
rect 13587 4505 13596 4539
rect 13544 4496 13596 4505
rect 7472 4428 7524 4480
rect 9956 4471 10008 4480
rect 9956 4437 9965 4471
rect 9965 4437 9999 4471
rect 9999 4437 10008 4471
rect 9956 4428 10008 4437
rect 15108 4496 15160 4548
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 16672 4607 16724 4616
rect 16672 4573 16681 4607
rect 16681 4573 16715 4607
rect 16715 4573 16724 4607
rect 16672 4564 16724 4573
rect 19340 4632 19392 4684
rect 20720 4632 20772 4684
rect 18696 4564 18748 4616
rect 19156 4564 19208 4616
rect 16948 4539 17000 4548
rect 16948 4505 16957 4539
rect 16957 4505 16991 4539
rect 16991 4505 17000 4539
rect 16948 4496 17000 4505
rect 15476 4428 15528 4480
rect 19340 4496 19392 4548
rect 22008 4607 22060 4616
rect 22008 4573 22017 4607
rect 22017 4573 22051 4607
rect 22051 4573 22060 4607
rect 22008 4564 22060 4573
rect 4266 4326 4318 4378
rect 4330 4326 4382 4378
rect 4394 4326 4446 4378
rect 4458 4326 4510 4378
rect 4522 4326 4574 4378
rect 9579 4326 9631 4378
rect 9643 4326 9695 4378
rect 9707 4326 9759 4378
rect 9771 4326 9823 4378
rect 9835 4326 9887 4378
rect 14892 4326 14944 4378
rect 14956 4326 15008 4378
rect 15020 4326 15072 4378
rect 15084 4326 15136 4378
rect 15148 4326 15200 4378
rect 20205 4326 20257 4378
rect 20269 4326 20321 4378
rect 20333 4326 20385 4378
rect 20397 4326 20449 4378
rect 20461 4326 20513 4378
rect 3976 4224 4028 4276
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 9956 4224 10008 4276
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 13544 4224 13596 4276
rect 13820 4224 13872 4276
rect 19064 4224 19116 4276
rect 4804 4156 4856 4208
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 5632 4156 5684 4208
rect 6276 4156 6328 4208
rect 17224 4156 17276 4208
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 7012 4088 7064 4140
rect 9404 4088 9456 4140
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 6920 4020 6972 4072
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 7380 4063 7432 4072
rect 7380 4029 7389 4063
rect 7389 4029 7423 4063
rect 7423 4029 7432 4063
rect 7380 4020 7432 4029
rect 7288 3952 7340 4004
rect 7656 3952 7708 4004
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 13544 4131 13596 4140
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 14004 4088 14056 4140
rect 13636 4063 13688 4072
rect 10784 3952 10836 4004
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 15476 4088 15528 4140
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 7748 3884 7800 3936
rect 11060 3884 11112 3936
rect 14004 3952 14056 4004
rect 16396 4020 16448 4072
rect 16672 4020 16724 4072
rect 19432 4156 19484 4208
rect 14556 3952 14608 4004
rect 19248 4063 19300 4072
rect 19248 4029 19257 4063
rect 19257 4029 19291 4063
rect 19291 4029 19300 4063
rect 19248 4020 19300 4029
rect 19340 4020 19392 4072
rect 19984 4020 20036 4072
rect 14096 3884 14148 3936
rect 16580 3884 16632 3936
rect 3606 3782 3658 3834
rect 3670 3782 3722 3834
rect 3734 3782 3786 3834
rect 3798 3782 3850 3834
rect 3862 3782 3914 3834
rect 8919 3782 8971 3834
rect 8983 3782 9035 3834
rect 9047 3782 9099 3834
rect 9111 3782 9163 3834
rect 9175 3782 9227 3834
rect 14232 3782 14284 3834
rect 14296 3782 14348 3834
rect 14360 3782 14412 3834
rect 14424 3782 14476 3834
rect 14488 3782 14540 3834
rect 19545 3782 19597 3834
rect 19609 3782 19661 3834
rect 19673 3782 19725 3834
rect 19737 3782 19789 3834
rect 19801 3782 19853 3834
rect 4896 3680 4948 3732
rect 6828 3680 6880 3732
rect 7380 3723 7432 3732
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 11980 3680 12032 3732
rect 13820 3680 13872 3732
rect 14004 3680 14056 3732
rect 16948 3680 17000 3732
rect 17040 3723 17092 3732
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 19248 3680 19300 3732
rect 6920 3612 6972 3664
rect 848 3408 900 3460
rect 6276 3544 6328 3596
rect 7288 3544 7340 3596
rect 7564 3544 7616 3596
rect 10600 3544 10652 3596
rect 6920 3476 6972 3528
rect 11244 3476 11296 3528
rect 11888 3476 11940 3528
rect 6644 3408 6696 3460
rect 10048 3408 10100 3460
rect 13636 3476 13688 3528
rect 13544 3451 13596 3460
rect 13544 3417 13553 3451
rect 13553 3417 13587 3451
rect 13587 3417 13596 3451
rect 13544 3408 13596 3417
rect 14188 3519 14240 3528
rect 14188 3485 14222 3519
rect 14222 3485 14240 3519
rect 14188 3476 14240 3485
rect 14648 3408 14700 3460
rect 16120 3544 16172 3596
rect 16488 3544 16540 3596
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16856 3519 16908 3528
rect 16396 3476 16448 3485
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 17316 3476 17368 3528
rect 19432 3519 19484 3528
rect 19432 3485 19440 3519
rect 19440 3485 19484 3519
rect 19432 3476 19484 3485
rect 17040 3408 17092 3460
rect 9956 3340 10008 3392
rect 14280 3340 14332 3392
rect 15292 3340 15344 3392
rect 17868 3340 17920 3392
rect 4266 3238 4318 3290
rect 4330 3238 4382 3290
rect 4394 3238 4446 3290
rect 4458 3238 4510 3290
rect 4522 3238 4574 3290
rect 9579 3238 9631 3290
rect 9643 3238 9695 3290
rect 9707 3238 9759 3290
rect 9771 3238 9823 3290
rect 9835 3238 9887 3290
rect 14892 3238 14944 3290
rect 14956 3238 15008 3290
rect 15020 3238 15072 3290
rect 15084 3238 15136 3290
rect 15148 3238 15200 3290
rect 20205 3238 20257 3290
rect 20269 3238 20321 3290
rect 20333 3238 20385 3290
rect 20397 3238 20449 3290
rect 20461 3238 20513 3290
rect 6920 3136 6972 3188
rect 9956 3136 10008 3188
rect 13544 3136 13596 3188
rect 14280 3179 14332 3188
rect 14280 3145 14289 3179
rect 14289 3145 14323 3179
rect 14323 3145 14332 3179
rect 14280 3136 14332 3145
rect 14648 3179 14700 3188
rect 14648 3145 14657 3179
rect 14657 3145 14691 3179
rect 14691 3145 14700 3179
rect 14648 3136 14700 3145
rect 16488 3136 16540 3188
rect 16856 3136 16908 3188
rect 17868 3136 17920 3188
rect 5540 3068 5592 3120
rect 6920 3043 6972 3052
rect 6920 3009 6938 3043
rect 6938 3009 6972 3043
rect 6920 3000 6972 3009
rect 10048 3000 10100 3052
rect 13820 3000 13872 3052
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 15016 3043 15068 3052
rect 15016 3009 15025 3043
rect 15025 3009 15059 3043
rect 15059 3009 15068 3043
rect 15016 3000 15068 3009
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 15292 2975 15344 2984
rect 15292 2941 15301 2975
rect 15301 2941 15335 2975
rect 15335 2941 15344 2975
rect 15292 2932 15344 2941
rect 19340 3068 19392 3120
rect 17316 3000 17368 3052
rect 20076 3000 20128 3052
rect 20628 2932 20680 2984
rect 7012 2796 7064 2848
rect 14188 2796 14240 2848
rect 14924 2796 14976 2848
rect 3606 2694 3658 2746
rect 3670 2694 3722 2746
rect 3734 2694 3786 2746
rect 3798 2694 3850 2746
rect 3862 2694 3914 2746
rect 8919 2694 8971 2746
rect 8983 2694 9035 2746
rect 9047 2694 9099 2746
rect 9111 2694 9163 2746
rect 9175 2694 9227 2746
rect 14232 2694 14284 2746
rect 14296 2694 14348 2746
rect 14360 2694 14412 2746
rect 14424 2694 14476 2746
rect 14488 2694 14540 2746
rect 19545 2694 19597 2746
rect 19609 2694 19661 2746
rect 19673 2694 19725 2746
rect 19737 2694 19789 2746
rect 19801 2694 19853 2746
rect 4804 2635 4856 2644
rect 4804 2601 4813 2635
rect 4813 2601 4847 2635
rect 4847 2601 4856 2635
rect 4804 2592 4856 2601
rect 5540 2592 5592 2644
rect 6920 2592 6972 2644
rect 10048 2592 10100 2644
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 11520 2592 11572 2644
rect 12532 2635 12584 2644
rect 12532 2601 12541 2635
rect 12541 2601 12575 2635
rect 12575 2601 12584 2635
rect 12532 2592 12584 2601
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 17040 2592 17092 2644
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 20076 2635 20128 2644
rect 20076 2601 20085 2635
rect 20085 2601 20119 2635
rect 20119 2601 20128 2635
rect 20076 2592 20128 2601
rect 3240 2388 3292 2440
rect 3884 2388 3936 2440
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5172 2388 5224 2440
rect 6460 2388 6512 2440
rect 7012 2456 7064 2508
rect 7288 2499 7340 2508
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 5816 2252 5868 2304
rect 6644 2295 6696 2304
rect 6644 2261 6653 2295
rect 6653 2261 6687 2295
rect 6687 2261 6696 2295
rect 6644 2252 6696 2261
rect 6920 2320 6972 2372
rect 7288 2320 7340 2372
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8576 2388 8628 2440
rect 9036 2388 9088 2440
rect 11336 2524 11388 2576
rect 12072 2524 12124 2576
rect 13820 2524 13872 2576
rect 15016 2524 15068 2576
rect 9956 2388 10008 2440
rect 10324 2388 10376 2440
rect 10968 2388 11020 2440
rect 11612 2388 11664 2440
rect 12256 2388 12308 2440
rect 13084 2388 13136 2440
rect 13544 2388 13596 2440
rect 13912 2388 13964 2440
rect 14740 2388 14792 2440
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 15568 2388 15620 2397
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 16764 2388 16816 2440
rect 17408 2388 17460 2440
rect 18052 2388 18104 2440
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 19340 2388 19392 2440
rect 19984 2388 20036 2440
rect 7196 2252 7248 2304
rect 7748 2252 7800 2304
rect 8392 2252 8444 2304
rect 11796 2320 11848 2372
rect 12900 2320 12952 2372
rect 11152 2252 11204 2304
rect 14188 2252 14240 2304
rect 15476 2252 15528 2304
rect 16120 2252 16172 2304
rect 16764 2252 16816 2304
rect 18696 2252 18748 2304
rect 4266 2150 4318 2202
rect 4330 2150 4382 2202
rect 4394 2150 4446 2202
rect 4458 2150 4510 2202
rect 4522 2150 4574 2202
rect 9579 2150 9631 2202
rect 9643 2150 9695 2202
rect 9707 2150 9759 2202
rect 9771 2150 9823 2202
rect 9835 2150 9887 2202
rect 14892 2150 14944 2202
rect 14956 2150 15008 2202
rect 15020 2150 15072 2202
rect 15084 2150 15136 2202
rect 15148 2150 15200 2202
rect 20205 2150 20257 2202
rect 20269 2150 20321 2202
rect 20333 2150 20385 2202
rect 20397 2150 20449 2202
rect 20461 2150 20513 2202
<< metal2 >>
rect 4526 24970 4582 25612
rect 5170 24970 5226 25612
rect 6458 24970 6514 25612
rect 4526 24942 4844 24970
rect 4526 24812 4582 24942
rect 3606 23420 3914 23429
rect 3606 23418 3612 23420
rect 3668 23418 3692 23420
rect 3748 23418 3772 23420
rect 3828 23418 3852 23420
rect 3908 23418 3914 23420
rect 3668 23366 3670 23418
rect 3850 23366 3852 23418
rect 3606 23364 3612 23366
rect 3668 23364 3692 23366
rect 3748 23364 3772 23366
rect 3828 23364 3852 23366
rect 3908 23364 3914 23366
rect 3606 23355 3914 23364
rect 4816 23118 4844 24942
rect 5170 24942 5304 24970
rect 5170 24812 5226 24942
rect 5276 23118 5304 24942
rect 6458 24942 6592 24970
rect 6458 24812 6514 24942
rect 6564 23118 6592 24942
rect 7102 24812 7158 25612
rect 7746 24970 7802 25612
rect 7746 24942 8064 24970
rect 7746 24812 7802 24942
rect 7116 23322 7144 24812
rect 8036 23322 8064 24942
rect 8390 24812 8446 25612
rect 9034 24970 9090 25612
rect 9034 24942 9352 24970
rect 9034 24812 9090 24942
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 8024 23316 8076 23322
rect 8024 23258 8076 23264
rect 8404 23118 8432 24812
rect 8919 23420 9227 23429
rect 8919 23418 8925 23420
rect 8981 23418 9005 23420
rect 9061 23418 9085 23420
rect 9141 23418 9165 23420
rect 9221 23418 9227 23420
rect 8981 23366 8983 23418
rect 9163 23366 9165 23418
rect 8919 23364 8925 23366
rect 8981 23364 9005 23366
rect 9061 23364 9085 23366
rect 9141 23364 9165 23366
rect 9221 23364 9227 23366
rect 8919 23355 9227 23364
rect 9324 23118 9352 24942
rect 9678 24812 9734 25612
rect 10322 24970 10378 25612
rect 10322 24942 10456 24970
rect 10322 24812 10378 24942
rect 9692 23118 9720 24812
rect 10428 23118 10456 24942
rect 10966 24812 11022 25612
rect 11610 24812 11666 25612
rect 12254 24812 12310 25612
rect 12898 24812 12954 25612
rect 13542 24812 13598 25612
rect 14186 24970 14242 25612
rect 14108 24942 14242 24970
rect 10980 23118 11008 24812
rect 11624 23322 11652 24812
rect 11612 23316 11664 23322
rect 11612 23258 11664 23264
rect 12268 23254 12296 24812
rect 11060 23248 11112 23254
rect 11060 23190 11112 23196
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 4804 23112 4856 23118
rect 4804 23054 4856 23060
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 10416 23112 10468 23118
rect 10416 23054 10468 23060
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 7288 23044 7340 23050
rect 7288 22986 7340 22992
rect 7932 23044 7984 23050
rect 7932 22986 7984 22992
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 4266 22876 4574 22885
rect 4266 22874 4272 22876
rect 4328 22874 4352 22876
rect 4408 22874 4432 22876
rect 4488 22874 4512 22876
rect 4568 22874 4574 22876
rect 4328 22822 4330 22874
rect 4510 22822 4512 22874
rect 4266 22820 4272 22822
rect 4328 22820 4352 22822
rect 4408 22820 4432 22822
rect 4488 22820 4512 22822
rect 4568 22820 4574 22822
rect 4266 22811 4574 22820
rect 846 22672 902 22681
rect 846 22607 848 22616
rect 900 22607 902 22616
rect 848 22578 900 22584
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 848 22024 900 22030
rect 846 21992 848 22001
rect 900 21992 902 22001
rect 846 21927 902 21936
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 848 21548 900 21554
rect 848 21490 900 21496
rect 860 21321 888 21490
rect 846 21312 902 21321
rect 846 21247 902 21256
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20505 1532 20742
rect 1490 20496 1546 20505
rect 1490 20431 1546 20440
rect 848 19712 900 19718
rect 846 19680 848 19689
rect 900 19680 902 19689
rect 846 19615 902 19624
rect 1492 19168 1544 19174
rect 1490 19136 1492 19145
rect 1544 19136 1546 19145
rect 1490 19071 1546 19080
rect 848 18760 900 18766
rect 848 18702 900 18708
rect 860 18601 888 18702
rect 846 18592 902 18601
rect 846 18527 902 18536
rect 1596 18426 1624 21830
rect 2700 21078 2728 22510
rect 3606 22332 3914 22341
rect 3606 22330 3612 22332
rect 3668 22330 3692 22332
rect 3748 22330 3772 22332
rect 3828 22330 3852 22332
rect 3908 22330 3914 22332
rect 3668 22278 3670 22330
rect 3850 22278 3852 22330
rect 3606 22276 3612 22278
rect 3668 22276 3692 22278
rect 3748 22276 3772 22278
rect 3828 22276 3852 22278
rect 3908 22276 3914 22278
rect 3606 22267 3914 22276
rect 4266 21788 4574 21797
rect 4266 21786 4272 21788
rect 4328 21786 4352 21788
rect 4408 21786 4432 21788
rect 4488 21786 4512 21788
rect 4568 21786 4574 21788
rect 4328 21734 4330 21786
rect 4510 21734 4512 21786
rect 4266 21732 4272 21734
rect 4328 21732 4352 21734
rect 4408 21732 4432 21734
rect 4488 21732 4512 21734
rect 4568 21732 4574 21734
rect 4266 21723 4574 21732
rect 4632 21554 4660 22918
rect 4896 22500 4948 22506
rect 4896 22442 4948 22448
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 3606 21244 3914 21253
rect 3606 21242 3612 21244
rect 3668 21242 3692 21244
rect 3748 21242 3772 21244
rect 3828 21242 3852 21244
rect 3908 21242 3914 21244
rect 3668 21190 3670 21242
rect 3850 21190 3852 21242
rect 3606 21188 3612 21190
rect 3668 21188 3692 21190
rect 3748 21188 3772 21190
rect 3828 21188 3852 21190
rect 3908 21188 3914 21190
rect 3606 21179 3914 21188
rect 2688 21072 2740 21078
rect 2688 21014 2740 21020
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1872 18290 1900 18566
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17785 1532 18022
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 848 17060 900 17066
rect 848 17002 900 17008
rect 860 16969 888 17002
rect 846 16960 902 16969
rect 846 16895 902 16904
rect 848 16584 900 16590
rect 846 16552 848 16561
rect 900 16552 902 16561
rect 846 16487 902 16496
rect 848 15904 900 15910
rect 846 15872 848 15881
rect 900 15872 902 15881
rect 846 15807 902 15816
rect 1780 15570 1808 17682
rect 1872 17678 1900 18226
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17746 1992 18022
rect 2424 17882 2452 18158
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 2516 17542 2544 18770
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2608 17678 2636 18362
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 2056 15434 2084 16390
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2424 15706 2452 16050
rect 2608 15706 2636 16050
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 2044 15428 2096 15434
rect 2044 15370 2096 15376
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1964 15162 1992 15302
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1398 15056 1454 15065
rect 2056 15026 2084 15370
rect 2148 15366 2176 15506
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 1398 14991 1454 15000
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2424 14958 2452 15642
rect 2608 15026 2636 15642
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 1676 14544 1728 14550
rect 846 14512 902 14521
rect 1676 14486 1728 14492
rect 846 14447 902 14456
rect 860 14414 888 14447
rect 848 14408 900 14414
rect 848 14350 900 14356
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 14074 1624 14214
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1688 13870 1716 14486
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 13161 888 13262
rect 846 13152 902 13161
rect 846 13087 902 13096
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 846 11792 902 11801
rect 846 11727 848 11736
rect 900 11727 902 11736
rect 1676 11756 1728 11762
rect 848 11698 900 11704
rect 1676 11698 1728 11704
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 10305 1532 11086
rect 1688 10985 1716 11698
rect 1780 11014 1808 11698
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1768 11008 1820 11014
rect 1674 10976 1730 10985
rect 1768 10950 1820 10956
rect 1674 10911 1730 10920
rect 1490 10296 1546 10305
rect 1490 10231 1546 10240
rect 1780 10062 1808 10950
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9625 1532 9862
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 848 9104 900 9110
rect 846 9072 848 9081
rect 900 9072 902 9081
rect 846 9007 902 9016
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8498 1716 8774
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1964 7954 1992 11018
rect 2240 10130 2268 11494
rect 2700 11286 2728 21014
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3988 20466 4016 20742
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3606 20156 3914 20165
rect 3606 20154 3612 20156
rect 3668 20154 3692 20156
rect 3748 20154 3772 20156
rect 3828 20154 3852 20156
rect 3908 20154 3914 20156
rect 3668 20102 3670 20154
rect 3850 20102 3852 20154
rect 3606 20100 3612 20102
rect 3668 20100 3692 20102
rect 3748 20100 3772 20102
rect 3828 20100 3852 20102
rect 3908 20100 3914 20102
rect 3606 20091 3914 20100
rect 4172 19310 4200 21422
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4540 21010 4568 21286
rect 4528 21004 4580 21010
rect 4528 20946 4580 20952
rect 4632 20874 4660 21490
rect 4908 21078 4936 22442
rect 5460 21690 5488 22918
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 4988 21412 5040 21418
rect 4988 21354 5040 21360
rect 4896 21072 4948 21078
rect 4896 21014 4948 21020
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4724 20874 4752 20946
rect 4908 20942 4936 21014
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 4266 20700 4574 20709
rect 4266 20698 4272 20700
rect 4328 20698 4352 20700
rect 4408 20698 4432 20700
rect 4488 20698 4512 20700
rect 4568 20698 4574 20700
rect 4328 20646 4330 20698
rect 4510 20646 4512 20698
rect 4266 20644 4272 20646
rect 4328 20644 4352 20646
rect 4408 20644 4432 20646
rect 4488 20644 4512 20646
rect 4568 20644 4574 20646
rect 4266 20635 4574 20644
rect 4266 19612 4574 19621
rect 4266 19610 4272 19612
rect 4328 19610 4352 19612
rect 4408 19610 4432 19612
rect 4488 19610 4512 19612
rect 4568 19610 4574 19612
rect 4328 19558 4330 19610
rect 4510 19558 4512 19610
rect 4266 19556 4272 19558
rect 4328 19556 4352 19558
rect 4408 19556 4432 19558
rect 4488 19556 4512 19558
rect 4568 19556 4574 19558
rect 4266 19547 4574 19556
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2792 18426 2820 18566
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2884 18290 2912 19246
rect 3606 19068 3914 19077
rect 3606 19066 3612 19068
rect 3668 19066 3692 19068
rect 3748 19066 3772 19068
rect 3828 19066 3852 19068
rect 3908 19066 3914 19068
rect 3668 19014 3670 19066
rect 3850 19014 3852 19066
rect 3606 19012 3612 19014
rect 3668 19012 3692 19014
rect 3748 19012 3772 19014
rect 3828 19012 3852 19014
rect 3908 19012 3914 19014
rect 3606 19003 3914 19012
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2884 16046 2912 18226
rect 2976 18154 3004 18702
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 18426 3372 18566
rect 4266 18524 4574 18533
rect 4266 18522 4272 18524
rect 4328 18522 4352 18524
rect 4408 18522 4432 18524
rect 4488 18522 4512 18524
rect 4568 18522 4574 18524
rect 4328 18470 4330 18522
rect 4510 18470 4512 18522
rect 4266 18468 4272 18470
rect 4328 18468 4352 18470
rect 4408 18468 4432 18470
rect 4488 18468 4512 18470
rect 4568 18468 4574 18470
rect 4266 18459 4574 18468
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2976 17814 3004 18090
rect 3606 17980 3914 17989
rect 3606 17978 3612 17980
rect 3668 17978 3692 17980
rect 3748 17978 3772 17980
rect 3828 17978 3852 17980
rect 3908 17978 3914 17980
rect 3668 17926 3670 17978
rect 3850 17926 3852 17978
rect 3606 17924 3612 17926
rect 3668 17924 3692 17926
rect 3748 17924 3772 17926
rect 3828 17924 3852 17926
rect 3908 17924 3914 17926
rect 3606 17915 3914 17924
rect 2964 17808 3016 17814
rect 2964 17750 3016 17756
rect 3988 17678 4016 18158
rect 4080 17814 4108 18226
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3606 16892 3914 16901
rect 3606 16890 3612 16892
rect 3668 16890 3692 16892
rect 3748 16890 3772 16892
rect 3828 16890 3852 16892
rect 3908 16890 3914 16892
rect 3668 16838 3670 16890
rect 3850 16838 3852 16890
rect 3606 16836 3612 16838
rect 3668 16836 3692 16838
rect 3748 16836 3772 16838
rect 3828 16836 3852 16838
rect 3908 16836 3914 16838
rect 3606 16827 3914 16836
rect 3988 16250 4016 17614
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2884 15638 2912 15982
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2884 12782 2912 15302
rect 3436 15162 3464 16050
rect 4172 16046 4200 18022
rect 4724 17882 4752 20810
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4816 19922 4844 20198
rect 5000 19938 5028 21354
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5552 20874 5580 21286
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5724 20868 5776 20874
rect 5724 20810 5776 20816
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5460 20602 5488 20742
rect 5448 20596 5500 20602
rect 5448 20538 5500 20544
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5368 19990 5396 20402
rect 5552 20262 5580 20810
rect 5736 20482 5764 20810
rect 5644 20454 5764 20482
rect 6000 20460 6052 20466
rect 5644 20398 5672 20454
rect 6000 20402 6052 20408
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4908 19910 5028 19938
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 4816 19310 4844 19858
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4816 18358 4844 18634
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 4908 18290 4936 19910
rect 5552 19854 5580 20198
rect 5644 19922 5672 20334
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5000 19378 5028 19790
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 5000 18970 5028 19314
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4908 17746 4936 18022
rect 5184 17746 5212 18702
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5644 18426 5672 18566
rect 5736 18426 5764 20198
rect 6012 20058 6040 20402
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 4266 17436 4574 17445
rect 4266 17434 4272 17436
rect 4328 17434 4352 17436
rect 4408 17434 4432 17436
rect 4488 17434 4512 17436
rect 4568 17434 4574 17436
rect 4328 17382 4330 17434
rect 4510 17382 4512 17434
rect 4266 17380 4272 17382
rect 4328 17380 4352 17382
rect 4408 17380 4432 17382
rect 4488 17380 4512 17382
rect 4568 17380 4574 17382
rect 4266 17371 4574 17380
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 4266 16348 4574 16357
rect 4266 16346 4272 16348
rect 4328 16346 4352 16348
rect 4408 16346 4432 16348
rect 4488 16346 4512 16348
rect 4568 16346 4574 16348
rect 4328 16294 4330 16346
rect 4510 16294 4512 16346
rect 4266 16292 4272 16294
rect 4328 16292 4352 16294
rect 4408 16292 4432 16294
rect 4488 16292 4512 16294
rect 4568 16292 4574 16294
rect 4266 16283 4574 16292
rect 5644 16250 5672 16526
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 3606 15804 3914 15813
rect 3606 15802 3612 15804
rect 3668 15802 3692 15804
rect 3748 15802 3772 15804
rect 3828 15802 3852 15804
rect 3908 15802 3914 15804
rect 3668 15750 3670 15802
rect 3850 15750 3852 15802
rect 3606 15748 3612 15750
rect 3668 15748 3692 15750
rect 3748 15748 3772 15750
rect 3828 15748 3852 15750
rect 3908 15748 3914 15750
rect 3606 15739 3914 15748
rect 3988 15502 4016 15982
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 15570 4108 15846
rect 4172 15638 4200 15982
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 15162 4200 15302
rect 4266 15260 4574 15269
rect 4266 15258 4272 15260
rect 4328 15258 4352 15260
rect 4408 15258 4432 15260
rect 4488 15258 4512 15260
rect 4568 15258 4574 15260
rect 4328 15206 4330 15258
rect 4510 15206 4512 15258
rect 4266 15204 4272 15206
rect 4328 15204 4352 15206
rect 4408 15204 4432 15206
rect 4488 15204 4512 15206
rect 4568 15204 4574 15206
rect 4266 15195 4574 15204
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4632 15094 4660 16050
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 3606 14716 3914 14725
rect 3606 14714 3612 14716
rect 3668 14714 3692 14716
rect 3748 14714 3772 14716
rect 3828 14714 3852 14716
rect 3908 14714 3914 14716
rect 3668 14662 3670 14714
rect 3850 14662 3852 14714
rect 3606 14660 3612 14662
rect 3668 14660 3692 14662
rect 3748 14660 3772 14662
rect 3828 14660 3852 14662
rect 3908 14660 3914 14662
rect 3606 14651 3914 14660
rect 4266 14172 4574 14181
rect 4266 14170 4272 14172
rect 4328 14170 4352 14172
rect 4408 14170 4432 14172
rect 4488 14170 4512 14172
rect 4568 14170 4574 14172
rect 4328 14118 4330 14170
rect 4510 14118 4512 14170
rect 4266 14116 4272 14118
rect 4328 14116 4352 14118
rect 4408 14116 4432 14118
rect 4488 14116 4512 14118
rect 4568 14116 4574 14118
rect 4266 14107 4574 14116
rect 4724 13938 4752 14894
rect 5368 14414 5396 15982
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15570 5488 15846
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5644 14958 5672 16050
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5736 14362 5764 18226
rect 5828 18222 5856 19178
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5920 18766 5948 19110
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5828 17746 5856 18158
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 5828 15638 5856 17682
rect 6012 17678 6040 18090
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6196 17202 6224 18022
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6196 15978 6224 17138
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 5908 15904 5960 15910
rect 5908 15846 5960 15852
rect 5920 15706 5948 15846
rect 6104 15706 6132 15914
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 5828 14482 5856 15574
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 6092 14408 6144 14414
rect 5368 13938 5396 14350
rect 5736 14334 5856 14362
rect 6092 14350 6144 14356
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 3606 13628 3914 13637
rect 3606 13626 3612 13628
rect 3668 13626 3692 13628
rect 3748 13626 3772 13628
rect 3828 13626 3852 13628
rect 3908 13626 3914 13628
rect 3668 13574 3670 13626
rect 3850 13574 3852 13626
rect 3606 13572 3612 13574
rect 3668 13572 3692 13574
rect 3748 13572 3772 13574
rect 3828 13572 3852 13574
rect 3908 13572 3914 13574
rect 3606 13563 3914 13572
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4172 12986 4200 13126
rect 4266 13084 4574 13093
rect 4266 13082 4272 13084
rect 4328 13082 4352 13084
rect 4408 13082 4432 13084
rect 4488 13082 4512 13084
rect 4568 13082 4574 13084
rect 4328 13030 4330 13082
rect 4510 13030 4512 13082
rect 4266 13028 4272 13030
rect 4328 13028 4352 13030
rect 4408 13028 4432 13030
rect 4488 13028 4512 13030
rect 4568 13028 4574 13030
rect 4266 13019 4574 13028
rect 4632 12986 4660 13194
rect 4908 12986 4936 13874
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 10266 2360 10542
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2148 9722 2176 10066
rect 2424 10062 2452 10678
rect 2976 10606 3004 10950
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 3068 10538 3096 11018
rect 3160 10674 3188 12650
rect 3606 12540 3914 12549
rect 3606 12538 3612 12540
rect 3668 12538 3692 12540
rect 3748 12538 3772 12540
rect 3828 12538 3852 12540
rect 3908 12538 3914 12540
rect 3668 12486 3670 12538
rect 3850 12486 3852 12538
rect 3606 12484 3612 12486
rect 3668 12484 3692 12486
rect 3748 12484 3772 12486
rect 3828 12484 3852 12486
rect 3908 12484 3914 12486
rect 3606 12475 3914 12484
rect 4172 12238 4200 12922
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4264 12442 4292 12718
rect 4632 12442 4660 12718
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4724 12238 4752 12854
rect 5092 12714 5120 13330
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4266 11996 4574 12005
rect 4266 11994 4272 11996
rect 4328 11994 4352 11996
rect 4408 11994 4432 11996
rect 4488 11994 4512 11996
rect 4568 11994 4574 11996
rect 4328 11942 4330 11994
rect 4510 11942 4512 11994
rect 4266 11940 4272 11942
rect 4328 11940 4352 11942
rect 4408 11940 4432 11942
rect 4488 11940 4512 11942
rect 4568 11940 4574 11942
rect 4266 11931 4574 11940
rect 3606 11452 3914 11461
rect 3606 11450 3612 11452
rect 3668 11450 3692 11452
rect 3748 11450 3772 11452
rect 3828 11450 3852 11452
rect 3908 11450 3914 11452
rect 3668 11398 3670 11450
rect 3850 11398 3852 11450
rect 3606 11396 3612 11398
rect 3668 11396 3692 11398
rect 3748 11396 3772 11398
rect 3828 11396 3852 11398
rect 3908 11396 3914 11398
rect 3606 11387 3914 11396
rect 5276 11218 5304 13874
rect 5368 13530 5396 13874
rect 5736 13530 5764 14214
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3252 10810 3280 10950
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3344 10674 3372 11086
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 3344 10470 3372 10610
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10198 3372 10406
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 3436 10130 3464 10542
rect 3606 10364 3914 10373
rect 3606 10362 3612 10364
rect 3668 10362 3692 10364
rect 3748 10362 3772 10364
rect 3828 10362 3852 10364
rect 3908 10362 3914 10364
rect 3668 10310 3670 10362
rect 3850 10310 3852 10362
rect 3606 10308 3612 10310
rect 3668 10308 3692 10310
rect 3748 10308 3772 10310
rect 3828 10308 3852 10310
rect 3908 10308 3914 10310
rect 3606 10299 3914 10308
rect 3988 10266 4016 11018
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10606 4108 10950
rect 4266 10908 4574 10917
rect 4266 10906 4272 10908
rect 4328 10906 4352 10908
rect 4408 10906 4432 10908
rect 4488 10906 4512 10908
rect 4568 10906 4574 10908
rect 4328 10854 4330 10906
rect 4510 10854 4512 10906
rect 4266 10852 4272 10854
rect 4328 10852 4352 10854
rect 4408 10852 4432 10854
rect 4488 10852 4512 10854
rect 4568 10852 4574 10854
rect 4266 10843 4574 10852
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4172 10198 4200 10406
rect 4540 10266 4568 10610
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1780 7546 1808 7686
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 846 7440 902 7449
rect 1872 7410 1900 7686
rect 846 7375 848 7384
rect 900 7375 902 7384
rect 1676 7404 1728 7410
rect 848 7346 900 7352
rect 1676 7346 1728 7352
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1688 6905 1716 7346
rect 1872 7274 1900 7346
rect 1964 7274 1992 7890
rect 2424 7478 2452 9998
rect 4172 9586 4200 10134
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4266 9820 4574 9829
rect 4266 9818 4272 9820
rect 4328 9818 4352 9820
rect 4408 9818 4432 9820
rect 4488 9818 4512 9820
rect 4568 9818 4574 9820
rect 4328 9766 4330 9818
rect 4510 9766 4512 9818
rect 4266 9764 4272 9766
rect 4328 9764 4352 9766
rect 4408 9764 4432 9766
rect 4488 9764 4512 9766
rect 4568 9764 4574 9766
rect 4266 9755 4574 9764
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4632 9518 4660 9998
rect 4724 9654 4752 11018
rect 5092 10810 5120 11086
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10130 4936 10406
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 5000 10062 5028 10474
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 3606 9276 3914 9285
rect 3606 9274 3612 9276
rect 3668 9274 3692 9276
rect 3748 9274 3772 9276
rect 3828 9274 3852 9276
rect 3908 9274 3914 9276
rect 3668 9222 3670 9274
rect 3850 9222 3852 9274
rect 3606 9220 3612 9222
rect 3668 9220 3692 9222
rect 3748 9220 3772 9222
rect 3828 9220 3852 9222
rect 3908 9220 3914 9222
rect 3606 9211 3914 9220
rect 4172 8634 4200 9386
rect 4266 8732 4574 8741
rect 4266 8730 4272 8732
rect 4328 8730 4352 8732
rect 4408 8730 4432 8732
rect 4488 8730 4512 8732
rect 4568 8730 4574 8732
rect 4328 8678 4330 8730
rect 4510 8678 4512 8730
rect 4266 8676 4272 8678
rect 4328 8676 4352 8678
rect 4408 8676 4432 8678
rect 4488 8676 4512 8678
rect 4568 8676 4574 8678
rect 4266 8667 4574 8676
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3068 8090 3096 8434
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2608 7546 2636 7686
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2412 7472 2464 7478
rect 2700 7426 2728 7686
rect 2412 7414 2464 7420
rect 2608 7410 2728 7426
rect 2596 7404 2728 7410
rect 2648 7398 2728 7404
rect 2596 7346 2648 7352
rect 1860 7268 1912 7274
rect 1860 7210 1912 7216
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 1674 6896 1730 6905
rect 1674 6831 1730 6840
rect 2608 6458 2636 7346
rect 3068 7342 3096 8026
rect 3252 7954 3280 8298
rect 3606 8188 3914 8197
rect 3606 8186 3612 8188
rect 3668 8186 3692 8188
rect 3748 8186 3772 8188
rect 3828 8186 3852 8188
rect 3908 8186 3914 8188
rect 3668 8134 3670 8186
rect 3850 8134 3852 8186
rect 3606 8132 3612 8134
rect 3668 8132 3692 8134
rect 3748 8132 3772 8134
rect 3828 8132 3852 8134
rect 3908 8132 3914 8134
rect 3606 8123 3914 8132
rect 4080 8090 4108 8434
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3252 7410 3280 7890
rect 4172 7478 4200 8434
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 7886 4292 8298
rect 4356 7954 4384 8502
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4266 7644 4574 7653
rect 4266 7642 4272 7644
rect 4328 7642 4352 7644
rect 4408 7642 4432 7644
rect 4488 7642 4512 7644
rect 4568 7642 4574 7644
rect 4328 7590 4330 7642
rect 4510 7590 4512 7642
rect 4266 7588 4272 7590
rect 4328 7588 4352 7590
rect 4408 7588 4432 7590
rect 4488 7588 4512 7590
rect 4568 7588 4574 7590
rect 4266 7579 4574 7588
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 3606 7100 3914 7109
rect 3606 7098 3612 7100
rect 3668 7098 3692 7100
rect 3748 7098 3772 7100
rect 3828 7098 3852 7100
rect 3908 7098 3914 7100
rect 3668 7046 3670 7098
rect 3850 7046 3852 7098
rect 3606 7044 3612 7046
rect 3668 7044 3692 7046
rect 3748 7044 3772 7046
rect 3828 7044 3852 7046
rect 3908 7044 3914 7046
rect 3606 7035 3914 7044
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 3344 5710 3372 6598
rect 4172 6440 4200 7210
rect 4266 6556 4574 6565
rect 4266 6554 4272 6556
rect 4328 6554 4352 6556
rect 4408 6554 4432 6556
rect 4488 6554 4512 6556
rect 4568 6554 4574 6556
rect 4328 6502 4330 6554
rect 4510 6502 4512 6554
rect 4266 6500 4272 6502
rect 4328 6500 4352 6502
rect 4408 6500 4432 6502
rect 4488 6500 4512 6502
rect 4568 6500 4574 6502
rect 4266 6491 4574 6500
rect 4172 6412 4292 6440
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 3528 5370 3556 6258
rect 3606 6012 3914 6021
rect 3606 6010 3612 6012
rect 3668 6010 3692 6012
rect 3748 6010 3772 6012
rect 3828 6010 3852 6012
rect 3908 6010 3914 6012
rect 3668 5958 3670 6010
rect 3850 5958 3852 6010
rect 3606 5956 3612 5958
rect 3668 5956 3692 5958
rect 3748 5956 3772 5958
rect 3828 5956 3852 5958
rect 3908 5956 3914 5958
rect 3606 5947 3914 5956
rect 3988 5914 4016 6258
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4080 5710 4108 6054
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5001 888 5170
rect 3988 5166 4016 5646
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5370 4108 5510
rect 4172 5370 4200 6258
rect 4264 5778 4292 6412
rect 4632 5794 4660 7754
rect 4724 7410 4752 8366
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4816 7342 4844 8434
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5092 7478 5120 7686
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4816 6458 4844 7278
rect 5276 6866 5304 11154
rect 5828 10742 5856 14334
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5920 13802 5948 13874
rect 6104 13870 6132 14350
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 13462 5948 13738
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6012 13274 6040 13330
rect 5920 13258 6040 13274
rect 5908 13252 6040 13258
rect 5960 13246 6040 13252
rect 5908 13194 5960 13200
rect 5920 12850 5948 13194
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10266 5856 10406
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5828 9042 5856 10202
rect 6288 9994 6316 16118
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6472 15502 6500 15982
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6472 14618 6500 15438
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6564 14414 6592 18634
rect 6656 18290 6684 18838
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 6748 16182 6776 16458
rect 6840 16250 6868 20946
rect 7024 20942 7052 22510
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7116 22166 7144 22374
rect 7104 22160 7156 22166
rect 7104 22102 7156 22108
rect 7116 21554 7144 22102
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7208 21010 7236 21286
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7208 20398 7236 20946
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7300 20244 7328 22986
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 22778 7788 22918
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7760 21978 7788 22034
rect 7760 21950 7880 21978
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7208 20216 7328 20244
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6932 17882 6960 18294
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7024 16454 7052 19722
rect 7208 18426 7236 20216
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19514 7328 19654
rect 7392 19514 7420 21830
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7484 20466 7512 20878
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7852 20330 7880 21950
rect 7840 20324 7892 20330
rect 7840 20266 7892 20272
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7576 19854 7604 20198
rect 7852 19922 7880 20266
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7380 19508 7432 19514
rect 7380 19450 7432 19456
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7392 18290 7420 19110
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7392 17882 7420 18226
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7484 16454 7512 19382
rect 7852 19242 7880 19858
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7852 18970 7880 19178
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7576 18290 7604 18566
rect 7944 18426 7972 22986
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 8404 22642 8432 22918
rect 9579 22876 9887 22885
rect 9579 22874 9585 22876
rect 9641 22874 9665 22876
rect 9721 22874 9745 22876
rect 9801 22874 9825 22876
rect 9881 22874 9887 22876
rect 9641 22822 9643 22874
rect 9823 22822 9825 22874
rect 9579 22820 9585 22822
rect 9641 22820 9665 22822
rect 9721 22820 9745 22822
rect 9801 22820 9825 22822
rect 9881 22820 9887 22822
rect 9579 22811 9887 22820
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8312 21690 8340 22374
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 8404 21570 8432 22578
rect 8919 22332 9227 22341
rect 8919 22330 8925 22332
rect 8981 22330 9005 22332
rect 9061 22330 9085 22332
rect 9141 22330 9165 22332
rect 9221 22330 9227 22332
rect 8981 22278 8983 22330
rect 9163 22278 9165 22330
rect 8919 22276 8925 22278
rect 8981 22276 9005 22278
rect 9061 22276 9085 22278
rect 9141 22276 9165 22278
rect 9221 22276 9227 22278
rect 8919 22267 9227 22276
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8036 21554 8432 21570
rect 8496 21554 8524 21966
rect 8024 21548 8432 21554
rect 8076 21542 8432 21548
rect 8484 21548 8536 21554
rect 8024 21490 8076 21496
rect 8484 21490 8536 21496
rect 8588 21418 8616 22034
rect 9579 21788 9887 21797
rect 9579 21786 9585 21788
rect 9641 21786 9665 21788
rect 9721 21786 9745 21788
rect 9801 21786 9825 21788
rect 9881 21786 9887 21788
rect 9641 21734 9643 21786
rect 9823 21734 9825 21786
rect 9579 21732 9585 21734
rect 9641 21732 9665 21734
rect 9721 21732 9745 21734
rect 9801 21732 9825 21734
rect 9881 21732 9887 21734
rect 9579 21723 9887 21732
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8312 20942 8340 21286
rect 8919 21244 9227 21253
rect 8919 21242 8925 21244
rect 8981 21242 9005 21244
rect 9061 21242 9085 21244
rect 9141 21242 9165 21244
rect 9221 21242 9227 21244
rect 8981 21190 8983 21242
rect 9163 21190 9165 21242
rect 8919 21188 8925 21190
rect 8981 21188 9005 21190
rect 9061 21188 9085 21190
rect 9141 21188 9165 21190
rect 9221 21188 9227 21190
rect 8919 21179 9227 21188
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9324 20466 9352 20742
rect 9579 20700 9887 20709
rect 9579 20698 9585 20700
rect 9641 20698 9665 20700
rect 9721 20698 9745 20700
rect 9801 20698 9825 20700
rect 9881 20698 9887 20700
rect 9641 20646 9643 20698
rect 9823 20646 9825 20698
rect 9579 20644 9585 20646
rect 9641 20644 9665 20646
rect 9721 20644 9745 20646
rect 9801 20644 9825 20646
rect 9881 20644 9887 20646
rect 9579 20635 9887 20644
rect 9968 20602 9996 22918
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 9312 20460 9364 20466
rect 9312 20402 9364 20408
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 8919 20156 9227 20165
rect 8919 20154 8925 20156
rect 8981 20154 9005 20156
rect 9061 20154 9085 20156
rect 9141 20154 9165 20156
rect 9221 20154 9227 20156
rect 8981 20102 8983 20154
rect 9163 20102 9165 20154
rect 8919 20100 8925 20102
rect 8981 20100 9005 20102
rect 9061 20100 9085 20102
rect 9141 20100 9165 20102
rect 9221 20100 9227 20102
rect 8919 20091 9227 20100
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 8772 19514 8800 19858
rect 9324 19854 9352 20402
rect 9416 19922 9444 20402
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 9579 19612 9887 19621
rect 9579 19610 9585 19612
rect 9641 19610 9665 19612
rect 9721 19610 9745 19612
rect 9801 19610 9825 19612
rect 9881 19610 9887 19612
rect 9641 19558 9643 19610
rect 9823 19558 9825 19610
rect 9579 19556 9585 19558
rect 9641 19556 9665 19558
rect 9721 19556 9745 19558
rect 9801 19556 9825 19558
rect 9881 19556 9887 19558
rect 9579 19547 9887 19556
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 18834 8432 19110
rect 8588 18834 8616 19314
rect 10060 19310 10088 19790
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 8919 19068 9227 19077
rect 8919 19066 8925 19068
rect 8981 19066 9005 19068
rect 9061 19066 9085 19068
rect 9141 19066 9165 19068
rect 9221 19066 9227 19068
rect 8981 19014 8983 19066
rect 9163 19014 9165 19066
rect 8919 19012 8925 19014
rect 8981 19012 9005 19014
rect 9061 19012 9085 19014
rect 9141 19012 9165 19014
rect 9221 19012 9227 19014
rect 8919 19003 9227 19012
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7576 17678 7604 18226
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7760 16590 7788 17546
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16658 8340 16934
rect 8496 16726 8524 17070
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 15026 7512 15846
rect 7760 15706 7788 16526
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8496 15450 8524 16662
rect 8588 16658 8616 18770
rect 9784 18766 9812 19110
rect 10152 18970 10180 19450
rect 10244 19242 10272 19858
rect 10428 19786 10456 20198
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10244 18766 10272 19178
rect 10428 18834 10456 19722
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 9579 18524 9887 18533
rect 9579 18522 9585 18524
rect 9641 18522 9665 18524
rect 9721 18522 9745 18524
rect 9801 18522 9825 18524
rect 9881 18522 9887 18524
rect 9641 18470 9643 18522
rect 9823 18470 9825 18522
rect 9579 18468 9585 18470
rect 9641 18468 9665 18470
rect 9721 18468 9745 18470
rect 9801 18468 9825 18470
rect 9881 18468 9887 18470
rect 9579 18459 9887 18468
rect 8919 17980 9227 17989
rect 8919 17978 8925 17980
rect 8981 17978 9005 17980
rect 9061 17978 9085 17980
rect 9141 17978 9165 17980
rect 9221 17978 9227 17980
rect 8981 17926 8983 17978
rect 9163 17926 9165 17978
rect 8919 17924 8925 17926
rect 8981 17924 9005 17926
rect 9061 17924 9085 17926
rect 9141 17924 9165 17926
rect 9221 17924 9227 17926
rect 8919 17915 9227 17924
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8588 15638 8616 16594
rect 8680 16114 8708 17478
rect 8864 17338 8892 17682
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8956 17338 8984 17614
rect 10152 17610 10180 17682
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 9579 17436 9887 17445
rect 9579 17434 9585 17436
rect 9641 17434 9665 17436
rect 9721 17434 9745 17436
rect 9801 17434 9825 17436
rect 9881 17434 9887 17436
rect 9641 17382 9643 17434
rect 9823 17382 9825 17434
rect 9579 17380 9585 17382
rect 9641 17380 9665 17382
rect 9721 17380 9745 17382
rect 9801 17380 9825 17382
rect 9881 17380 9887 17382
rect 9579 17371 9887 17380
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 10152 17134 10180 17546
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10520 17134 10548 17206
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 8919 16892 9227 16901
rect 8919 16890 8925 16892
rect 8981 16890 9005 16892
rect 9061 16890 9085 16892
rect 9141 16890 9165 16892
rect 9221 16890 9227 16892
rect 8981 16838 8983 16890
rect 9163 16838 9165 16890
rect 8919 16836 8925 16838
rect 8981 16836 9005 16838
rect 9061 16836 9085 16838
rect 9141 16836 9165 16838
rect 9221 16836 9227 16838
rect 8919 16827 9227 16836
rect 10520 16658 10548 17070
rect 10704 16794 10732 20266
rect 10796 19446 10824 20334
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10520 16454 10548 16594
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 9579 16348 9887 16357
rect 9579 16346 9585 16348
rect 9641 16346 9665 16348
rect 9721 16346 9745 16348
rect 9801 16346 9825 16348
rect 9881 16346 9887 16348
rect 9641 16294 9643 16346
rect 9823 16294 9825 16346
rect 9579 16292 9585 16294
rect 9641 16292 9665 16294
rect 9721 16292 9745 16294
rect 9801 16292 9825 16294
rect 9881 16292 9887 16294
rect 9579 16283 9887 16292
rect 10520 16250 10548 16390
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 8919 15804 9227 15813
rect 8919 15802 8925 15804
rect 8981 15802 9005 15804
rect 9061 15802 9085 15804
rect 9141 15802 9165 15804
rect 9221 15802 9227 15804
rect 8981 15750 8983 15802
rect 9163 15750 9165 15802
rect 8919 15748 8925 15750
rect 8981 15748 9005 15750
rect 9061 15748 9085 15750
rect 9141 15748 9165 15750
rect 9221 15748 9227 15750
rect 8919 15739 9227 15748
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 10520 15570 10548 15846
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 8312 15422 8524 15450
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 7760 15162 7788 15370
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13870 6408 14214
rect 8128 13870 8156 14962
rect 8312 14958 8340 15422
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 14482 8340 14894
rect 8496 14890 8524 15302
rect 8588 15162 8616 15438
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 9579 15260 9887 15269
rect 9579 15258 9585 15260
rect 9641 15258 9665 15260
rect 9721 15258 9745 15260
rect 9801 15258 9825 15260
rect 9881 15258 9887 15260
rect 9641 15206 9643 15258
rect 9823 15206 9825 15258
rect 9579 15204 9585 15206
rect 9641 15204 9665 15206
rect 9721 15204 9745 15206
rect 9801 15204 9825 15206
rect 9881 15204 9887 15206
rect 9579 15195 9887 15204
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8772 14618 8800 14894
rect 8919 14716 9227 14725
rect 8919 14714 8925 14716
rect 8981 14714 9005 14716
rect 9061 14714 9085 14716
rect 9141 14714 9165 14716
rect 9221 14714 9227 14716
rect 8981 14662 8983 14714
rect 9163 14662 9165 14714
rect 8919 14660 8925 14662
rect 8981 14660 9005 14662
rect 9061 14660 9085 14662
rect 9141 14660 9165 14662
rect 9221 14660 9227 14662
rect 8919 14651 9227 14660
rect 9416 14618 9444 14962
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 9220 14408 9272 14414
rect 9272 14368 9352 14396
rect 9220 14350 9272 14356
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 13938 8708 14214
rect 9324 14074 9352 14368
rect 9508 14346 9536 14554
rect 9680 14544 9732 14550
rect 9864 14544 9916 14550
rect 9732 14492 9864 14498
rect 9680 14486 9916 14492
rect 9692 14470 9904 14486
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8220 13530 8248 13874
rect 9324 13870 9352 14010
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 8919 13628 9227 13637
rect 8919 13626 8925 13628
rect 8981 13626 9005 13628
rect 9061 13626 9085 13628
rect 9141 13626 9165 13628
rect 9221 13626 9227 13628
rect 8981 13574 8983 13626
rect 9163 13574 9165 13626
rect 8919 13572 8925 13574
rect 8981 13572 9005 13574
rect 9061 13572 9085 13574
rect 9141 13572 9165 13574
rect 9221 13572 9227 13574
rect 8919 13563 9227 13572
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 9324 13394 9352 13806
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12374 6960 12582
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6932 12186 6960 12310
rect 6932 12158 7144 12186
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6932 11898 6960 12038
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7024 11762 7052 12038
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 7546 5396 7686
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5460 7426 5488 7958
rect 5552 7886 5580 8298
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 7954 5672 8230
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5368 7398 5488 7426
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 4712 6248 4764 6254
rect 4764 6196 4936 6202
rect 4712 6190 4936 6196
rect 4724 6186 4936 6190
rect 4724 6180 4948 6186
rect 4724 6174 4896 6180
rect 4896 6122 4948 6128
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4252 5772 4304 5778
rect 4632 5766 4752 5794
rect 4252 5714 4304 5720
rect 4264 5574 4292 5714
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4266 5468 4574 5477
rect 4266 5466 4272 5468
rect 4328 5466 4352 5468
rect 4408 5466 4432 5468
rect 4488 5466 4512 5468
rect 4568 5466 4574 5468
rect 4328 5414 4330 5466
rect 4510 5414 4512 5466
rect 4266 5412 4272 5414
rect 4328 5412 4352 5414
rect 4408 5412 4432 5414
rect 4488 5412 4512 5414
rect 4568 5412 4574 5414
rect 4266 5403 4574 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4632 5302 4660 5646
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 846 4992 902 5001
rect 846 4927 902 4936
rect 3606 4924 3914 4933
rect 3606 4922 3612 4924
rect 3668 4922 3692 4924
rect 3748 4922 3772 4924
rect 3828 4922 3852 4924
rect 3908 4922 3914 4924
rect 3668 4870 3670 4922
rect 3850 4870 3852 4922
rect 3606 4868 3612 4870
rect 3668 4868 3692 4870
rect 3748 4868 3772 4870
rect 3828 4868 3852 4870
rect 3908 4868 3914 4870
rect 3606 4859 3914 4868
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 860 4321 888 4558
rect 846 4312 902 4321
rect 3988 4282 4016 5102
rect 4724 4690 4752 5766
rect 4816 5370 4844 6054
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 5000 5302 5028 6326
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 5092 4826 5120 6666
rect 5276 6458 5304 6666
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5368 6254 5396 7398
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5460 6390 5488 6734
rect 5552 6662 5580 7686
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6012 6866 6040 7278
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6104 6458 6132 6598
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 6104 5914 6132 6258
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5460 5234 5488 5714
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5736 5166 5764 5646
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4266 4380 4574 4389
rect 4266 4378 4272 4380
rect 4328 4378 4352 4380
rect 4408 4378 4432 4380
rect 4488 4378 4512 4380
rect 4568 4378 4574 4380
rect 4328 4326 4330 4378
rect 4510 4326 4512 4378
rect 4266 4324 4272 4326
rect 4328 4324 4352 4326
rect 4408 4324 4432 4326
rect 4488 4324 4512 4326
rect 4568 4324 4574 4326
rect 4266 4315 4574 4324
rect 846 4247 902 4256
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 4724 4078 4752 4626
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5644 4214 5672 4558
rect 6288 4214 6316 9930
rect 6380 8974 6408 11494
rect 7024 11218 7052 11698
rect 7116 11558 7144 12158
rect 7208 11694 7236 12786
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 7116 11150 7144 11494
rect 7300 11218 7328 11630
rect 7392 11626 7420 12038
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7288 11212 7340 11218
rect 7340 11172 7420 11200
rect 7288 11154 7340 11160
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6748 10674 6776 11018
rect 7208 10674 7236 11154
rect 7392 10742 7420 11172
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9178 6500 9862
rect 6748 9586 6776 9998
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6748 9178 6776 9522
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6840 7886 6868 9522
rect 6932 8838 6960 9998
rect 7208 9586 7236 10066
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7300 8974 7328 10406
rect 7392 9042 7420 10678
rect 7576 10538 7604 12718
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7668 12306 7696 12650
rect 8919 12540 9227 12549
rect 8919 12538 8925 12540
rect 8981 12538 9005 12540
rect 9061 12538 9085 12540
rect 9141 12538 9165 12540
rect 9221 12538 9227 12540
rect 8981 12486 8983 12538
rect 9163 12486 9165 12538
rect 8919 12484 8925 12486
rect 8981 12484 9005 12486
rect 9061 12484 9085 12486
rect 9141 12484 9165 12486
rect 9221 12484 9227 12486
rect 8919 12475 9227 12484
rect 9416 12442 9444 14214
rect 9508 14056 9536 14282
rect 9579 14172 9887 14181
rect 9579 14170 9585 14172
rect 9641 14170 9665 14172
rect 9721 14170 9745 14172
rect 9801 14170 9825 14172
rect 9881 14170 9887 14172
rect 9641 14118 9643 14170
rect 9823 14118 9825 14170
rect 9579 14116 9585 14118
rect 9641 14116 9665 14118
rect 9721 14116 9745 14118
rect 9801 14116 9825 14118
rect 9881 14116 9887 14118
rect 9579 14107 9887 14116
rect 9508 14028 9720 14056
rect 9692 13938 9720 14028
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9692 13462 9720 13874
rect 9968 13870 9996 14350
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 10060 13802 10088 13942
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 10060 13258 10088 13738
rect 10152 13326 10180 14554
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10244 14074 10272 14486
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10336 13394 10364 13670
rect 10520 13394 10548 15370
rect 10612 15366 10640 15982
rect 10704 15434 10732 16730
rect 10796 16522 10824 17002
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10796 15706 10824 16458
rect 10888 16114 10916 22918
rect 10980 22574 11008 22918
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 20398 11008 22510
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 11072 19718 11100 23190
rect 12912 23118 12940 24812
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 12808 23044 12860 23050
rect 12808 22986 12860 22992
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11072 19378 11100 19654
rect 11164 19514 11192 19654
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 11256 19446 11284 19654
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10980 17746 11008 19110
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11164 17338 11192 17546
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11716 16114 11744 22918
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10888 15502 10916 16050
rect 11900 15706 11928 22986
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 21962 12480 22374
rect 12636 22166 12664 22918
rect 12624 22160 12676 22166
rect 12624 22102 12676 22108
rect 12636 21962 12664 22102
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 12452 21486 12480 21898
rect 12636 21554 12664 21898
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12636 21418 12664 21490
rect 12624 21412 12676 21418
rect 12624 21354 12676 21360
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12544 18698 12572 19858
rect 12728 19854 12756 21830
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12820 19514 12848 22986
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13096 22778 13124 22918
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 13372 22574 13400 23122
rect 13556 23118 13584 24812
rect 14108 23322 14136 24942
rect 14186 24812 14242 24942
rect 14830 24970 14886 25612
rect 15474 24970 15530 25612
rect 14830 24942 15148 24970
rect 14830 24812 14886 24942
rect 14232 23420 14540 23429
rect 14232 23418 14238 23420
rect 14294 23418 14318 23420
rect 14374 23418 14398 23420
rect 14454 23418 14478 23420
rect 14534 23418 14540 23420
rect 14294 23366 14296 23418
rect 14476 23366 14478 23418
rect 14232 23364 14238 23366
rect 14294 23364 14318 23366
rect 14374 23364 14398 23366
rect 14454 23364 14478 23366
rect 14534 23364 14540 23366
rect 14232 23355 14540 23364
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 15120 23118 15148 24942
rect 15474 24942 15608 24970
rect 15474 24812 15530 24942
rect 15580 23118 15608 24942
rect 16118 24812 16174 25612
rect 16762 24812 16818 25612
rect 17406 24812 17462 25612
rect 18050 24970 18106 25612
rect 18694 24970 18750 25612
rect 19338 24970 19394 25612
rect 18050 24942 18368 24970
rect 18050 24812 18106 24942
rect 16132 23254 16160 24812
rect 16776 23322 16804 24812
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16120 23248 16172 23254
rect 16120 23190 16172 23196
rect 17420 23118 17448 24812
rect 18340 23322 18368 24942
rect 18694 24942 19012 24970
rect 18694 24812 18750 24942
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18984 23118 19012 24942
rect 19338 24942 19472 24970
rect 19338 24812 19394 24942
rect 19444 23118 19472 24942
rect 19545 23420 19853 23429
rect 19545 23418 19551 23420
rect 19607 23418 19631 23420
rect 19687 23418 19711 23420
rect 19767 23418 19791 23420
rect 19847 23418 19853 23420
rect 19607 23366 19609 23418
rect 19789 23366 19791 23418
rect 19545 23364 19551 23366
rect 19607 23364 19631 23366
rect 19687 23364 19711 23366
rect 19767 23364 19791 23366
rect 19847 23364 19853 23366
rect 19545 23355 19853 23364
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13912 22976 13964 22982
rect 13912 22918 13964 22924
rect 13648 22642 13676 22918
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13924 22574 13952 22918
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13188 20466 13216 21286
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 13096 19378 13124 20334
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13188 19310 13216 20402
rect 13280 19922 13308 22034
rect 13372 20058 13400 22510
rect 13924 22098 13952 22510
rect 13912 22092 13964 22098
rect 13912 22034 13964 22040
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13740 21486 13768 21966
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 13464 20942 13492 21286
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13648 20534 13676 20810
rect 13636 20528 13688 20534
rect 13636 20470 13688 20476
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 13280 19310 13308 19654
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12544 17066 12572 18634
rect 13372 18408 13400 19994
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13188 18380 13400 18408
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 17678 12756 18090
rect 12912 17746 12940 18158
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 17270 12756 17614
rect 12912 17270 12940 17682
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12912 16726 12940 17206
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 13004 16794 13032 17070
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 13188 16658 13216 18380
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16250 12572 16390
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12636 16046 12664 16594
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10612 13870 10640 15302
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 11532 13394 11560 13942
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11808 13326 11836 13874
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 9579 13084 9887 13093
rect 9579 13082 9585 13084
rect 9641 13082 9665 13084
rect 9721 13082 9745 13084
rect 9801 13082 9825 13084
rect 9881 13082 9887 13084
rect 9641 13030 9643 13082
rect 9823 13030 9825 13082
rect 9579 13028 9585 13030
rect 9641 13028 9665 13030
rect 9721 13028 9745 13030
rect 9801 13028 9825 13030
rect 9881 13028 9887 13030
rect 9579 13019 9887 13028
rect 12084 12986 12112 13126
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12176 12458 12204 15914
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12360 13394 12388 13942
rect 12452 13870 12480 14350
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12636 13530 12664 13874
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12268 12850 12296 13126
rect 12360 12918 12388 13330
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 13190 12848 13262
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 9404 12436 9456 12442
rect 12176 12430 12388 12458
rect 12544 12442 12572 12718
rect 9404 12378 9456 12384
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8036 11626 8064 11698
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11150 7696 11494
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 8128 11082 8156 12242
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 8944 12164 8996 12170
rect 8944 12106 8996 12112
rect 8956 11898 8984 12106
rect 9579 11996 9887 12005
rect 9579 11994 9585 11996
rect 9641 11994 9665 11996
rect 9721 11994 9745 11996
rect 9801 11994 9825 11996
rect 9881 11994 9887 11996
rect 9641 11942 9643 11994
rect 9823 11942 9825 11994
rect 9579 11940 9585 11942
rect 9641 11940 9665 11942
rect 9721 11940 9745 11942
rect 9801 11940 9825 11942
rect 9881 11940 9887 11942
rect 9579 11931 9887 11940
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 10152 11694 10180 12174
rect 10428 11762 10456 12242
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10428 11626 10456 11698
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 8588 11354 8616 11562
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 8919 11452 9227 11461
rect 8919 11450 8925 11452
rect 8981 11450 9005 11452
rect 9061 11450 9085 11452
rect 9141 11450 9165 11452
rect 9221 11450 9227 11452
rect 8981 11398 8983 11450
rect 9163 11398 9165 11450
rect 8919 11396 8925 11398
rect 8981 11396 9005 11398
rect 9061 11396 9085 11398
rect 9141 11396 9165 11398
rect 9221 11396 9227 11398
rect 8919 11387 9227 11396
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 9416 11150 9444 11494
rect 10428 11354 10456 11562
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7852 10742 7880 11018
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7576 9722 7604 10474
rect 8128 10266 8156 11018
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 9048 10810 9076 10950
rect 9579 10908 9887 10917
rect 9579 10906 9585 10908
rect 9641 10906 9665 10908
rect 9721 10906 9745 10908
rect 9801 10906 9825 10908
rect 9881 10906 9887 10908
rect 9641 10854 9643 10906
rect 9823 10854 9825 10906
rect 9579 10852 9585 10854
rect 9641 10852 9665 10854
rect 9721 10852 9745 10854
rect 9801 10852 9825 10854
rect 9881 10852 9887 10854
rect 9579 10843 9887 10852
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 10244 10742 10272 10950
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7760 8974 7788 9522
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 8220 8498 8248 10406
rect 8919 10364 9227 10373
rect 8919 10362 8925 10364
rect 8981 10362 9005 10364
rect 9061 10362 9085 10364
rect 9141 10362 9165 10364
rect 9221 10362 9227 10364
rect 8981 10310 8983 10362
rect 9163 10310 9165 10362
rect 8919 10308 8925 10310
rect 8981 10308 9005 10310
rect 9061 10308 9085 10310
rect 9141 10308 9165 10310
rect 9221 10308 9227 10310
rect 8919 10299 9227 10308
rect 8919 9276 9227 9285
rect 8919 9274 8925 9276
rect 8981 9274 9005 9276
rect 9061 9274 9085 9276
rect 9141 9274 9165 9276
rect 9221 9274 9227 9276
rect 8981 9222 8983 9274
rect 9163 9222 9165 9274
rect 8919 9220 8925 9222
rect 8981 9220 9005 9222
rect 9061 9220 9085 9222
rect 9141 9220 9165 9222
rect 9221 9220 9227 9222
rect 8919 9211 9227 9220
rect 9416 9110 9444 10542
rect 10428 10062 10456 11290
rect 10612 11150 10640 11494
rect 10980 11286 11008 11630
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10266 10732 10950
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10980 10062 11008 11222
rect 11348 11218 11376 11698
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11348 10742 11376 11154
rect 11808 11082 11836 11154
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11532 10690 11560 10950
rect 11624 10810 11652 10950
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11532 10674 11652 10690
rect 11532 10668 11664 10674
rect 11532 10662 11612 10668
rect 11612 10610 11664 10616
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 9579 9820 9887 9829
rect 9579 9818 9585 9820
rect 9641 9818 9665 9820
rect 9721 9818 9745 9820
rect 9801 9818 9825 9820
rect 9881 9818 9887 9820
rect 9641 9766 9643 9818
rect 9823 9766 9825 9818
rect 9579 9764 9585 9766
rect 9641 9764 9665 9766
rect 9721 9764 9745 9766
rect 9801 9764 9825 9766
rect 9881 9764 9887 9766
rect 9579 9755 9887 9764
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9416 8514 9444 9046
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9508 8634 9536 8842
rect 9579 8732 9887 8741
rect 9579 8730 9585 8732
rect 9641 8730 9665 8732
rect 9721 8730 9745 8732
rect 9801 8730 9825 8732
rect 9881 8730 9887 8732
rect 9641 8678 9643 8730
rect 9823 8678 9825 8730
rect 9579 8676 9585 8678
rect 9641 8676 9665 8678
rect 9721 8676 9745 8678
rect 9801 8676 9825 8678
rect 9881 8676 9887 8678
rect 9579 8667 9887 8676
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 10232 8560 10284 8566
rect 8208 8492 8260 8498
rect 9416 8486 9536 8514
rect 10232 8502 10284 8508
rect 8208 8434 8260 8440
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7002 6868 7822
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6564 6186 6592 6802
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6458 6868 6734
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 7024 5710 7052 6190
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 3606 3836 3914 3845
rect 3606 3834 3612 3836
rect 3668 3834 3692 3836
rect 3748 3834 3772 3836
rect 3828 3834 3852 3836
rect 3908 3834 3914 3836
rect 3668 3782 3670 3834
rect 3850 3782 3852 3834
rect 3606 3780 3612 3782
rect 3668 3780 3692 3782
rect 3748 3780 3772 3782
rect 3828 3780 3852 3782
rect 3908 3780 3914 3782
rect 3606 3771 3914 3780
rect 848 3460 900 3466
rect 848 3402 900 3408
rect 860 3369 888 3402
rect 846 3360 902 3369
rect 846 3295 902 3304
rect 4266 3292 4574 3301
rect 4266 3290 4272 3292
rect 4328 3290 4352 3292
rect 4408 3290 4432 3292
rect 4488 3290 4512 3292
rect 4568 3290 4574 3292
rect 4328 3238 4330 3290
rect 4510 3238 4512 3290
rect 4266 3236 4272 3238
rect 4328 3236 4352 3238
rect 4408 3236 4432 3238
rect 4488 3236 4512 3238
rect 4568 3236 4574 3238
rect 4266 3227 4574 3236
rect 3606 2748 3914 2757
rect 3606 2746 3612 2748
rect 3668 2746 3692 2748
rect 3748 2746 3772 2748
rect 3828 2746 3852 2748
rect 3908 2746 3914 2748
rect 3668 2694 3670 2746
rect 3850 2694 3852 2746
rect 3606 2692 3612 2694
rect 3668 2692 3692 2694
rect 3748 2692 3772 2694
rect 3828 2692 3852 2694
rect 3908 2692 3914 2694
rect 3606 2683 3914 2692
rect 4816 2650 4844 4150
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3738 4936 4082
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 6288 3602 6316 4150
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6656 3466 6684 4082
rect 6840 3738 6868 5170
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6932 4078 6960 4558
rect 7024 4146 7052 4626
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6932 3670 6960 4014
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6932 3534 6960 3606
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5552 2650 5580 3062
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 3252 800 3280 2382
rect 3896 800 3924 2382
rect 4266 2204 4574 2213
rect 4266 2202 4272 2204
rect 4328 2202 4352 2204
rect 4408 2202 4432 2204
rect 4488 2202 4512 2204
rect 4568 2202 4574 2204
rect 4328 2150 4330 2202
rect 4510 2150 4512 2202
rect 4266 2148 4272 2150
rect 4328 2148 4352 2150
rect 4408 2148 4432 2150
rect 4488 2148 4512 2150
rect 4568 2148 4574 2150
rect 4266 2139 4574 2148
rect 4632 1306 4660 2382
rect 4540 1278 4660 1306
rect 4540 800 4568 1278
rect 5184 800 5212 2382
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 800 5856 2246
rect 6472 800 6500 2382
rect 6656 2310 6684 3402
rect 6932 3194 6960 3470
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6932 2650 6960 2994
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6932 2378 6960 2586
rect 7024 2514 7052 2790
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7116 2394 7144 8298
rect 8220 7886 8248 8434
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 8919 8188 9227 8197
rect 8919 8186 8925 8188
rect 8981 8186 9005 8188
rect 9061 8186 9085 8188
rect 9141 8186 9165 8188
rect 9221 8186 9227 8188
rect 8981 8134 8983 8186
rect 9163 8134 9165 8186
rect 8919 8132 8925 8134
rect 8981 8132 9005 8134
rect 9061 8132 9085 8134
rect 9141 8132 9165 8134
rect 9221 8132 9227 8134
rect 8919 8123 9227 8132
rect 9324 8090 9352 8366
rect 9416 8294 9444 8366
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9416 7886 9444 8230
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 7208 7546 7236 7822
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7208 4078 7236 5646
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7300 4010 7328 5102
rect 7392 4162 7420 7686
rect 7668 7410 7696 7822
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7668 6458 7696 7346
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7576 5914 7604 6190
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4282 7512 4422
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7392 4134 7512 4162
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7392 3738 7420 4014
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7300 2514 7328 3538
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7484 2446 7512 4134
rect 7576 3602 7604 5510
rect 7668 4010 7696 6258
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7760 3942 7788 4490
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7760 2990 7788 3878
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7852 2446 7880 7142
rect 8404 6798 8432 7754
rect 8919 7100 9227 7109
rect 8919 7098 8925 7100
rect 8981 7098 9005 7100
rect 9061 7098 9085 7100
rect 9141 7098 9165 7100
rect 9221 7098 9227 7100
rect 8981 7046 8983 7098
rect 9163 7046 9165 7098
rect 8919 7044 8925 7046
rect 8981 7044 9005 7046
rect 9061 7044 9085 7046
rect 9141 7044 9165 7046
rect 9221 7044 9227 7046
rect 8919 7035 9227 7044
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8404 6458 8432 6734
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5914 8156 6054
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7944 5166 7972 5510
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 8588 2446 8616 6598
rect 9508 6440 9536 8486
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9600 8362 9628 8434
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9600 7954 9628 8298
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 9579 7644 9887 7653
rect 9579 7642 9585 7644
rect 9641 7642 9665 7644
rect 9721 7642 9745 7644
rect 9801 7642 9825 7644
rect 9881 7642 9887 7644
rect 9641 7590 9643 7642
rect 9823 7590 9825 7642
rect 9579 7588 9585 7590
rect 9641 7588 9665 7590
rect 9721 7588 9745 7590
rect 9801 7588 9825 7590
rect 9881 7588 9887 7590
rect 9579 7579 9887 7588
rect 9968 7478 9996 7686
rect 10152 7478 10180 7686
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 9579 6556 9887 6565
rect 9579 6554 9585 6556
rect 9641 6554 9665 6556
rect 9721 6554 9745 6556
rect 9801 6554 9825 6556
rect 9881 6554 9887 6556
rect 9641 6502 9643 6554
rect 9823 6502 9825 6554
rect 9579 6500 9585 6502
rect 9641 6500 9665 6502
rect 9721 6500 9745 6502
rect 9801 6500 9825 6502
rect 9881 6500 9887 6502
rect 9579 6491 9887 6500
rect 9416 6412 9536 6440
rect 9416 6254 9444 6412
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 8919 6012 9227 6021
rect 8919 6010 8925 6012
rect 8981 6010 9005 6012
rect 9061 6010 9085 6012
rect 9141 6010 9165 6012
rect 9221 6010 9227 6012
rect 8981 5958 8983 6010
rect 9163 5958 9165 6010
rect 8919 5956 8925 5958
rect 8981 5956 9005 5958
rect 9061 5956 9085 5958
rect 9141 5956 9165 5958
rect 9221 5956 9227 5958
rect 8919 5947 9227 5956
rect 8919 4924 9227 4933
rect 8919 4922 8925 4924
rect 8981 4922 9005 4924
rect 9061 4922 9085 4924
rect 9141 4922 9165 4924
rect 9221 4922 9227 4924
rect 8981 4870 8983 4922
rect 9163 4870 9165 4922
rect 8919 4868 8925 4870
rect 8981 4868 9005 4870
rect 9061 4868 9085 4870
rect 9141 4868 9165 4870
rect 9221 4868 9227 4870
rect 8919 4859 9227 4868
rect 9508 4758 9536 6258
rect 9784 5914 9812 6258
rect 10244 6254 10272 8502
rect 10336 7886 10364 8910
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 7886 10456 8774
rect 10612 8498 10640 8842
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10336 7290 10364 7822
rect 10336 7262 10456 7290
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 10244 5846 10272 6190
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10060 5642 10088 5714
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9579 5468 9887 5477
rect 9579 5466 9585 5468
rect 9641 5466 9665 5468
rect 9721 5466 9745 5468
rect 9801 5466 9825 5468
rect 9881 5466 9887 5468
rect 9641 5414 9643 5466
rect 9823 5414 9825 5466
rect 9579 5412 9585 5414
rect 9641 5412 9665 5414
rect 9721 5412 9745 5414
rect 9801 5412 9825 5414
rect 9881 5412 9887 5414
rect 9579 5403 9887 5412
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 4826 9628 5170
rect 10060 4826 10088 5578
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 10244 4690 10272 5782
rect 10336 5778 10364 7142
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 9416 4146 9444 4626
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9579 4380 9887 4389
rect 9579 4378 9585 4380
rect 9641 4378 9665 4380
rect 9721 4378 9745 4380
rect 9801 4378 9825 4380
rect 9881 4378 9887 4380
rect 9641 4326 9643 4378
rect 9823 4326 9825 4378
rect 9579 4324 9585 4326
rect 9641 4324 9665 4326
rect 9721 4324 9745 4326
rect 9801 4324 9825 4326
rect 9881 4324 9887 4326
rect 9579 4315 9887 4324
rect 9968 4282 9996 4422
rect 10152 4282 10180 4490
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 8919 3836 9227 3845
rect 8919 3834 8925 3836
rect 8981 3834 9005 3836
rect 9061 3834 9085 3836
rect 9141 3834 9165 3836
rect 9221 3834 9227 3836
rect 8981 3782 8983 3834
rect 9163 3782 9165 3834
rect 8919 3780 8925 3782
rect 8981 3780 9005 3782
rect 9061 3780 9085 3782
rect 9141 3780 9165 3782
rect 9221 3780 9227 3782
rect 8919 3771 9227 3780
rect 9416 3738 9444 4082
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9579 3292 9887 3301
rect 9579 3290 9585 3292
rect 9641 3290 9665 3292
rect 9721 3290 9745 3292
rect 9801 3290 9825 3292
rect 9881 3290 9887 3292
rect 9641 3238 9643 3290
rect 9823 3238 9825 3290
rect 9579 3236 9585 3238
rect 9641 3236 9665 3238
rect 9721 3236 9745 3238
rect 9801 3236 9825 3238
rect 9881 3236 9887 3238
rect 9579 3227 9887 3236
rect 9968 3194 9996 3334
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10060 3058 10088 3402
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 8919 2748 9227 2757
rect 8919 2746 8925 2748
rect 8981 2746 9005 2748
rect 9061 2746 9085 2748
rect 9141 2746 9165 2748
rect 9221 2746 9227 2748
rect 8981 2694 8983 2746
rect 9163 2694 9165 2746
rect 8919 2692 8925 2694
rect 8981 2692 9005 2694
rect 9061 2692 9085 2694
rect 9141 2692 9165 2694
rect 9221 2692 9227 2694
rect 8919 2683 9227 2692
rect 10060 2650 10088 2994
rect 10428 2650 10456 7262
rect 10612 3602 10640 7822
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10704 5302 10732 5850
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10796 4010 10824 4626
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 11072 3942 11100 8910
rect 11348 8514 11376 8910
rect 11532 8566 11560 8978
rect 11164 8486 11376 8514
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 7472 2440 7524 2446
rect 7116 2378 7328 2394
rect 7472 2382 7524 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 6920 2372 6972 2378
rect 7116 2372 7340 2378
rect 7116 2366 7288 2372
rect 6920 2314 6972 2320
rect 7288 2314 7340 2320
rect 6644 2304 6696 2310
rect 7196 2304 7248 2310
rect 6644 2246 6696 2252
rect 7116 2264 7196 2292
rect 7116 800 7144 2264
rect 7196 2246 7248 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 9048 800 9076 2382
rect 9579 2204 9887 2213
rect 9579 2202 9585 2204
rect 9641 2202 9665 2204
rect 9721 2202 9745 2204
rect 9801 2202 9825 2204
rect 9881 2202 9887 2204
rect 9641 2150 9643 2202
rect 9823 2150 9825 2202
rect 9579 2148 9585 2150
rect 9641 2148 9665 2150
rect 9721 2148 9745 2150
rect 9801 2148 9825 2150
rect 9881 2148 9887 2150
rect 9579 2139 9887 2148
rect 9692 870 9812 898
rect 9692 800 9720 870
rect 18 0 74 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 9784 762 9812 870
rect 9968 762 9996 2382
rect 10336 800 10364 2382
rect 10980 800 11008 2382
rect 11164 2310 11192 8486
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11256 7954 11284 8366
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11256 2650 11284 3470
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11348 2582 11376 7822
rect 11624 2774 11652 10610
rect 11808 5778 11836 11018
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10674 11928 10950
rect 12084 10810 12112 11018
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5370 11836 5510
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11900 5250 11928 10610
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11532 2746 11652 2774
rect 11808 5222 11928 5250
rect 11532 2650 11560 2746
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11624 800 11652 2382
rect 11808 2378 11836 5222
rect 11992 5166 12020 10406
rect 12360 10062 12388 12430
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12636 12238 12664 12786
rect 12820 12782 12848 13126
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 11218 12572 11494
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12912 10062 12940 14758
rect 13004 14074 13032 14962
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13096 14618 13124 14894
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13096 12986 13124 13194
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12268 8090 12296 8366
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12452 8022 12480 9862
rect 12728 9722 12756 9998
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12820 9654 12848 9998
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12544 8090 12572 8910
rect 12728 8566 12756 8910
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12360 6322 12388 7210
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12084 6186 12112 6258
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12084 5234 12112 5646
rect 12360 5370 12388 6258
rect 12544 6186 12572 7346
rect 12636 6866 12664 8434
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13004 7546 13032 7686
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 13096 7478 13124 7686
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13096 6322 13124 6802
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13188 6202 13216 10202
rect 13280 9994 13308 18090
rect 13372 17882 13400 18226
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13464 17814 13492 19858
rect 13832 19514 13860 19926
rect 14016 19514 14044 22986
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 14108 22098 14136 22646
rect 14232 22332 14540 22341
rect 14232 22330 14238 22332
rect 14294 22330 14318 22332
rect 14374 22330 14398 22332
rect 14454 22330 14478 22332
rect 14534 22330 14540 22332
rect 14294 22278 14296 22330
rect 14476 22278 14478 22330
rect 14232 22276 14238 22278
rect 14294 22276 14318 22278
rect 14374 22276 14398 22278
rect 14454 22276 14478 22278
rect 14534 22276 14540 22278
rect 14232 22267 14540 22276
rect 14096 22092 14148 22098
rect 14096 22034 14148 22040
rect 14232 21244 14540 21253
rect 14232 21242 14238 21244
rect 14294 21242 14318 21244
rect 14374 21242 14398 21244
rect 14454 21242 14478 21244
rect 14534 21242 14540 21244
rect 14294 21190 14296 21242
rect 14476 21190 14478 21242
rect 14232 21188 14238 21190
rect 14294 21188 14318 21190
rect 14374 21188 14398 21190
rect 14454 21188 14478 21190
rect 14534 21188 14540 21190
rect 14232 21179 14540 21188
rect 14232 20156 14540 20165
rect 14232 20154 14238 20156
rect 14294 20154 14318 20156
rect 14374 20154 14398 20156
rect 14454 20154 14478 20156
rect 14534 20154 14540 20156
rect 14294 20102 14296 20154
rect 14476 20102 14478 20154
rect 14232 20100 14238 20102
rect 14294 20100 14318 20102
rect 14374 20100 14398 20102
rect 14454 20100 14478 20102
rect 14534 20100 14540 20102
rect 14232 20091 14540 20100
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13556 18426 13584 19314
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13832 18358 13860 19450
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13924 18290 13952 19314
rect 14108 18902 14136 19790
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14476 19310 14504 19722
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14232 19068 14540 19077
rect 14232 19066 14238 19068
rect 14294 19066 14318 19068
rect 14374 19066 14398 19068
rect 14454 19066 14478 19068
rect 14534 19066 14540 19068
rect 14294 19014 14296 19066
rect 14476 19014 14478 19066
rect 14232 19012 14238 19014
rect 14294 19012 14318 19014
rect 14374 19012 14398 19014
rect 14454 19012 14478 19014
rect 14534 19012 14540 19014
rect 14232 19003 14540 19012
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14108 18358 14136 18838
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13464 17218 13492 17750
rect 13464 17190 13584 17218
rect 13556 17134 13584 17190
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13464 16114 13492 16526
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13556 16250 13584 16390
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13648 15502 13676 18226
rect 14232 17980 14540 17989
rect 14232 17978 14238 17980
rect 14294 17978 14318 17980
rect 14374 17978 14398 17980
rect 14454 17978 14478 17980
rect 14534 17978 14540 17980
rect 14294 17926 14296 17978
rect 14476 17926 14478 17978
rect 14232 17924 14238 17926
rect 14294 17924 14318 17926
rect 14374 17924 14398 17926
rect 14454 17924 14478 17926
rect 14534 17924 14540 17926
rect 14232 17915 14540 17924
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13648 15162 13676 15438
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14482 13584 14758
rect 13740 14482 13768 17070
rect 14232 16892 14540 16901
rect 14232 16890 14238 16892
rect 14294 16890 14318 16892
rect 14374 16890 14398 16892
rect 14454 16890 14478 16892
rect 14534 16890 14540 16892
rect 14294 16838 14296 16890
rect 14476 16838 14478 16890
rect 14232 16836 14238 16838
rect 14294 16836 14318 16838
rect 14374 16836 14398 16838
rect 14454 16836 14478 16838
rect 14534 16836 14540 16838
rect 14232 16827 14540 16836
rect 13820 16516 13872 16522
rect 13820 16458 13872 16464
rect 13832 16182 13860 16458
rect 14568 16182 14596 22918
rect 14892 22876 15200 22885
rect 14892 22874 14898 22876
rect 14954 22874 14978 22876
rect 15034 22874 15058 22876
rect 15114 22874 15138 22876
rect 15194 22874 15200 22876
rect 14954 22822 14956 22874
rect 15136 22822 15138 22874
rect 14892 22820 14898 22822
rect 14954 22820 14978 22822
rect 15034 22820 15058 22822
rect 15114 22820 15138 22822
rect 15194 22820 15200 22822
rect 14892 22811 15200 22820
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14660 19514 14688 21830
rect 14892 21788 15200 21797
rect 14892 21786 14898 21788
rect 14954 21786 14978 21788
rect 15034 21786 15058 21788
rect 15114 21786 15138 21788
rect 15194 21786 15200 21788
rect 14954 21734 14956 21786
rect 15136 21734 15138 21786
rect 14892 21732 14898 21734
rect 14954 21732 14978 21734
rect 15034 21732 15058 21734
rect 15114 21732 15138 21734
rect 15194 21732 15200 21734
rect 14892 21723 15200 21732
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14892 20700 15200 20709
rect 14892 20698 14898 20700
rect 14954 20698 14978 20700
rect 15034 20698 15058 20700
rect 15114 20698 15138 20700
rect 15194 20698 15200 20700
rect 14954 20646 14956 20698
rect 15136 20646 15138 20698
rect 14892 20644 14898 20646
rect 14954 20644 14978 20646
rect 15034 20644 15058 20646
rect 15114 20644 15138 20646
rect 15194 20644 15200 20646
rect 14892 20635 15200 20644
rect 15304 20466 15332 20878
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15212 19854 15240 20198
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19514 14780 19654
rect 14892 19612 15200 19621
rect 14892 19610 14898 19612
rect 14954 19610 14978 19612
rect 15034 19610 15058 19612
rect 15114 19610 15138 19612
rect 15194 19610 15200 19612
rect 14954 19558 14956 19610
rect 15136 19558 15138 19610
rect 14892 19556 14898 19558
rect 14954 19556 14978 19558
rect 15034 19556 15058 19558
rect 15114 19556 15138 19558
rect 15194 19556 15200 19558
rect 14892 19547 15200 19556
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14892 18524 15200 18533
rect 14892 18522 14898 18524
rect 14954 18522 14978 18524
rect 15034 18522 15058 18524
rect 15114 18522 15138 18524
rect 15194 18522 15200 18524
rect 14954 18470 14956 18522
rect 15136 18470 15138 18522
rect 14892 18468 14898 18470
rect 14954 18468 14978 18470
rect 15034 18468 15058 18470
rect 15114 18468 15138 18470
rect 15194 18468 15200 18470
rect 14892 18459 15200 18468
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 14892 17436 15200 17445
rect 14892 17434 14898 17436
rect 14954 17434 14978 17436
rect 15034 17434 15058 17436
rect 15114 17434 15138 17436
rect 15194 17434 15200 17436
rect 14954 17382 14956 17434
rect 15136 17382 15138 17434
rect 14892 17380 14898 17382
rect 14954 17380 14978 17382
rect 15034 17380 15058 17382
rect 15114 17380 15138 17382
rect 15194 17380 15200 17382
rect 14892 17371 15200 17380
rect 15304 17338 15332 17478
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15396 17218 15424 22918
rect 15672 22642 15700 23054
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 15752 22976 15804 22982
rect 15752 22918 15804 22924
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15488 22098 15516 22374
rect 15764 22166 15792 22918
rect 16132 22778 16160 22918
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 16500 22642 16528 22918
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16684 22438 16712 22578
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 15488 21622 15516 22034
rect 15476 21616 15528 21622
rect 15476 21558 15528 21564
rect 15488 21486 15516 21558
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15580 20058 15608 22034
rect 15672 21078 15700 22034
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 21690 15976 21830
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 16132 21554 16160 22034
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15660 21072 15712 21078
rect 15660 21014 15712 21020
rect 15672 20398 15700 21014
rect 15856 20874 15884 21286
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15660 20392 15712 20398
rect 16776 20346 16804 22986
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17144 20466 17172 20878
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 15660 20334 15712 20340
rect 16684 20318 16804 20346
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15304 17190 15424 17218
rect 15304 16590 15332 17190
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 14892 16348 15200 16357
rect 14892 16346 14898 16348
rect 14954 16346 14978 16348
rect 15034 16346 15058 16348
rect 15114 16346 15138 16348
rect 15194 16346 15200 16348
rect 14954 16294 14956 16346
rect 15136 16294 15138 16346
rect 14892 16292 14898 16294
rect 14954 16292 14978 16294
rect 15034 16292 15058 16294
rect 15114 16292 15138 16294
rect 15194 16292 15200 16294
rect 14892 16283 15200 16292
rect 15396 16250 15424 16458
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14232 15804 14540 15813
rect 14232 15802 14238 15804
rect 14294 15802 14318 15804
rect 14374 15802 14398 15804
rect 14454 15802 14478 15804
rect 14534 15802 14540 15804
rect 14294 15750 14296 15802
rect 14476 15750 14478 15802
rect 14232 15748 14238 15750
rect 14294 15748 14318 15750
rect 14374 15748 14398 15750
rect 14454 15748 14478 15750
rect 14534 15748 14540 15750
rect 14232 15739 14540 15748
rect 14892 15260 15200 15269
rect 14892 15258 14898 15260
rect 14954 15258 14978 15260
rect 15034 15258 15058 15260
rect 15114 15258 15138 15260
rect 15194 15258 15200 15260
rect 14954 15206 14956 15258
rect 15136 15206 15138 15258
rect 14892 15204 14898 15206
rect 14954 15204 14978 15206
rect 15034 15204 15058 15206
rect 15114 15204 15138 15206
rect 15194 15204 15200 15206
rect 14892 15195 15200 15204
rect 15488 15042 15516 19722
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15856 18290 15884 19450
rect 16684 18426 16712 20318
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 16776 19854 16804 20198
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 17052 19514 17080 20198
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17144 19514 17172 19654
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15764 16658 15792 17138
rect 15856 16794 15884 18226
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15396 15014 15516 15042
rect 14232 14716 14540 14725
rect 14232 14714 14238 14716
rect 14294 14714 14318 14716
rect 14374 14714 14398 14716
rect 14454 14714 14478 14716
rect 14534 14714 14540 14716
rect 14294 14662 14296 14714
rect 14476 14662 14478 14714
rect 14232 14660 14238 14662
rect 14294 14660 14318 14662
rect 14374 14660 14398 14662
rect 14454 14660 14478 14662
rect 14534 14660 14540 14662
rect 14232 14651 14540 14660
rect 15396 14618 15424 15014
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14618 15516 14894
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13372 13870 13400 14214
rect 13740 13938 13768 14214
rect 14660 14074 14688 14350
rect 14892 14172 15200 14181
rect 14892 14170 14898 14172
rect 14954 14170 14978 14172
rect 15034 14170 15058 14172
rect 15114 14170 15138 14172
rect 15194 14170 15200 14172
rect 14954 14118 14956 14170
rect 15136 14118 15138 14170
rect 14892 14116 14898 14118
rect 14954 14116 14978 14118
rect 15034 14116 15058 14118
rect 15114 14116 15138 14118
rect 15194 14116 15200 14118
rect 14892 14107 15200 14116
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13648 13326 13676 13806
rect 14232 13628 14540 13637
rect 14232 13626 14238 13628
rect 14294 13626 14318 13628
rect 14374 13626 14398 13628
rect 14454 13626 14478 13628
rect 14534 13626 14540 13628
rect 14294 13574 14296 13626
rect 14476 13574 14478 13626
rect 14232 13572 14238 13574
rect 14294 13572 14318 13574
rect 14374 13572 14398 13574
rect 14454 13572 14478 13574
rect 14534 13572 14540 13574
rect 14232 13563 14540 13572
rect 14660 13394 14688 14010
rect 15304 13870 15332 14486
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15396 13938 15424 14214
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15488 13870 15516 14554
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15304 13530 15332 13806
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13372 12918 13400 13194
rect 14892 13084 15200 13093
rect 14892 13082 14898 13084
rect 14954 13082 14978 13084
rect 15034 13082 15058 13084
rect 15114 13082 15138 13084
rect 15194 13082 15200 13084
rect 14954 13030 14956 13082
rect 15136 13030 15138 13082
rect 14892 13028 14898 13030
rect 14954 13028 14978 13030
rect 15034 13028 15058 13030
rect 15114 13028 15138 13030
rect 15194 13028 15200 13030
rect 14892 13019 15200 13028
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 14232 12540 14540 12549
rect 14232 12538 14238 12540
rect 14294 12538 14318 12540
rect 14374 12538 14398 12540
rect 14454 12538 14478 12540
rect 14534 12538 14540 12540
rect 14294 12486 14296 12538
rect 14476 12486 14478 12538
rect 14232 12484 14238 12486
rect 14294 12484 14318 12486
rect 14374 12484 14398 12486
rect 14454 12484 14478 12486
rect 14534 12484 14540 12486
rect 14232 12475 14540 12484
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13636 11212 13688 11218
rect 13832 11200 13860 11698
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14016 11218 14044 11630
rect 14108 11218 14136 12310
rect 14892 11996 15200 12005
rect 14892 11994 14898 11996
rect 14954 11994 14978 11996
rect 15034 11994 15058 11996
rect 15114 11994 15138 11996
rect 15194 11994 15200 11996
rect 14954 11942 14956 11994
rect 15136 11942 15138 11994
rect 14892 11940 14898 11942
rect 14954 11940 14978 11942
rect 15034 11940 15058 11942
rect 15114 11940 15138 11942
rect 15194 11940 15200 11942
rect 14892 11931 15200 11940
rect 15304 11762 15332 12582
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14232 11452 14540 11461
rect 14232 11450 14238 11452
rect 14294 11450 14318 11452
rect 14374 11450 14398 11452
rect 14454 11450 14478 11452
rect 14534 11450 14540 11452
rect 14294 11398 14296 11450
rect 14476 11398 14478 11450
rect 14232 11396 14238 11398
rect 14294 11396 14318 11398
rect 14374 11396 14398 11398
rect 14454 11396 14478 11398
rect 14534 11396 14540 11398
rect 14232 11387 14540 11396
rect 13688 11172 13860 11200
rect 13636 11154 13688 11160
rect 13832 10538 13860 11172
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14016 10606 14044 11154
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 14108 10470 14136 11154
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14476 10538 14504 10950
rect 14568 10606 14596 11494
rect 14752 10674 14780 11494
rect 15396 11286 15424 12650
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15200 11008 15252 11014
rect 15252 10968 15332 10996
rect 15200 10950 15252 10956
rect 14892 10908 15200 10917
rect 14892 10906 14898 10908
rect 14954 10906 14978 10908
rect 15034 10906 15058 10908
rect 15114 10906 15138 10908
rect 15194 10906 15200 10908
rect 14954 10854 14956 10906
rect 15136 10854 15138 10906
rect 14892 10852 14898 10854
rect 14954 10852 14978 10854
rect 15034 10852 15058 10854
rect 15114 10852 15138 10854
rect 15194 10852 15200 10854
rect 14892 10843 15200 10852
rect 15304 10742 15332 10968
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 14232 10364 14540 10373
rect 14232 10362 14238 10364
rect 14294 10362 14318 10364
rect 14374 10362 14398 10364
rect 14454 10362 14478 10364
rect 14534 10362 14540 10364
rect 14294 10310 14296 10362
rect 14476 10310 14478 10362
rect 14232 10308 14238 10310
rect 14294 10308 14318 10310
rect 14374 10308 14398 10310
rect 14454 10308 14478 10310
rect 14534 10308 14540 10310
rect 14232 10299 14540 10308
rect 14660 10062 14688 10406
rect 15304 10130 15332 10406
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 15396 9994 15424 10202
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14232 9276 14540 9285
rect 14232 9274 14238 9276
rect 14294 9274 14318 9276
rect 14374 9274 14398 9276
rect 14454 9274 14478 9276
rect 14534 9274 14540 9276
rect 14294 9222 14296 9274
rect 14476 9222 14478 9274
rect 14232 9220 14238 9222
rect 14294 9220 14318 9222
rect 14374 9220 14398 9222
rect 14454 9220 14478 9222
rect 14534 9220 14540 9222
rect 14232 9211 14540 9220
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13372 8498 13400 8910
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13280 7954 13308 8434
rect 14232 8188 14540 8197
rect 14232 8186 14238 8188
rect 14294 8186 14318 8188
rect 14374 8186 14398 8188
rect 14454 8186 14478 8188
rect 14534 8186 14540 8188
rect 14294 8134 14296 8186
rect 14476 8134 14478 8186
rect 14232 8132 14238 8134
rect 14294 8132 14318 8134
rect 14374 8132 14398 8134
rect 14454 8132 14478 8134
rect 14534 8132 14540 8134
rect 14232 8123 14540 8132
rect 14568 7954 14596 9862
rect 14660 8974 14688 9862
rect 14892 9820 15200 9829
rect 14892 9818 14898 9820
rect 14954 9818 14978 9820
rect 15034 9818 15058 9820
rect 15114 9818 15138 9820
rect 15194 9818 15200 9820
rect 14954 9766 14956 9818
rect 15136 9766 15138 9818
rect 14892 9764 14898 9766
rect 14954 9764 14978 9766
rect 15034 9764 15058 9766
rect 15114 9764 15138 9766
rect 15194 9764 15200 9766
rect 14892 9755 15200 9764
rect 15396 9654 15424 9930
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14752 8820 14780 9522
rect 15396 9110 15424 9590
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 14660 8792 14780 8820
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 13096 6174 13216 6202
rect 12544 5914 12572 6122
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 13004 5710 13032 6054
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11900 3534 11928 4082
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11992 3738 12020 4014
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 12084 2582 12112 5170
rect 12544 2650 12572 5578
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 13096 2446 13124 6174
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13188 5710 13216 6054
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13832 5574 13860 6258
rect 13924 6254 13952 6734
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13740 4622 13768 5102
rect 13832 4706 13860 5510
rect 13924 4826 13952 6190
rect 14016 5846 14044 7890
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14108 6186 14136 7346
rect 14232 7100 14540 7109
rect 14232 7098 14238 7100
rect 14294 7098 14318 7100
rect 14374 7098 14398 7100
rect 14454 7098 14478 7100
rect 14534 7098 14540 7100
rect 14294 7046 14296 7098
rect 14476 7046 14478 7098
rect 14232 7044 14238 7046
rect 14294 7044 14318 7046
rect 14374 7044 14398 7046
rect 14454 7044 14478 7046
rect 14534 7044 14540 7046
rect 14232 7035 14540 7044
rect 14660 6866 14688 8792
rect 14892 8732 15200 8741
rect 14892 8730 14898 8732
rect 14954 8730 14978 8732
rect 15034 8730 15058 8732
rect 15114 8730 15138 8732
rect 15194 8730 15200 8732
rect 14954 8678 14956 8730
rect 15136 8678 15138 8730
rect 14892 8676 14898 8678
rect 14954 8676 14978 8678
rect 15034 8676 15058 8678
rect 15114 8676 15138 8678
rect 15194 8676 15200 8678
rect 14892 8667 15200 8676
rect 15304 8498 15332 9046
rect 15488 8974 15516 10474
rect 15580 10198 15608 16390
rect 16316 16250 16344 16526
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15672 14618 15700 16050
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15844 16040 15896 16046
rect 16408 15994 16436 17682
rect 15844 15982 15896 15988
rect 15764 15706 15792 15982
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15856 15094 15884 15982
rect 16316 15978 16436 15994
rect 16304 15972 16436 15978
rect 16356 15966 16436 15972
rect 16304 15914 16356 15920
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15570 16252 15846
rect 16316 15570 16344 15914
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 16132 14958 16160 15302
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16316 14618 16344 15506
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16500 14618 16528 14962
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16028 14544 16080 14550
rect 16080 14492 16344 14498
rect 16028 14486 16344 14492
rect 16040 14482 16344 14486
rect 16040 14476 16356 14482
rect 16040 14470 16304 14476
rect 16304 14418 16356 14424
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 14074 16712 14214
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 17052 12238 17080 18294
rect 17328 18154 17356 22986
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17512 20398 17540 20878
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17880 20058 17908 20334
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17420 18222 17448 19246
rect 18064 18442 18092 22986
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 20942 19472 22918
rect 20205 22876 20513 22885
rect 20205 22874 20211 22876
rect 20267 22874 20291 22876
rect 20347 22874 20371 22876
rect 20427 22874 20451 22876
rect 20507 22874 20513 22876
rect 20267 22822 20269 22874
rect 20449 22822 20451 22874
rect 20205 22820 20211 22822
rect 20267 22820 20291 22822
rect 20347 22820 20371 22822
rect 20427 22820 20451 22822
rect 20507 22820 20513 22822
rect 20205 22811 20513 22820
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19545 22332 19853 22341
rect 19545 22330 19551 22332
rect 19607 22330 19631 22332
rect 19687 22330 19711 22332
rect 19767 22330 19791 22332
rect 19847 22330 19853 22332
rect 19607 22278 19609 22330
rect 19789 22278 19791 22330
rect 19545 22276 19551 22278
rect 19607 22276 19631 22278
rect 19687 22276 19711 22278
rect 19767 22276 19791 22278
rect 19847 22276 19853 22278
rect 19545 22267 19853 22276
rect 19545 21244 19853 21253
rect 19545 21242 19551 21244
rect 19607 21242 19631 21244
rect 19687 21242 19711 21244
rect 19767 21242 19791 21244
rect 19847 21242 19853 21244
rect 19607 21190 19609 21242
rect 19789 21190 19791 21242
rect 19545 21188 19551 21190
rect 19607 21188 19631 21190
rect 19687 21188 19711 21190
rect 19767 21188 19791 21190
rect 19847 21188 19853 21190
rect 19545 21179 19853 21188
rect 19904 21010 19932 22374
rect 20205 21788 20513 21797
rect 20205 21786 20211 21788
rect 20267 21786 20291 21788
rect 20347 21786 20371 21788
rect 20427 21786 20451 21788
rect 20507 21786 20513 21788
rect 20267 21734 20269 21786
rect 20449 21734 20451 21786
rect 20205 21732 20211 21734
rect 20267 21732 20291 21734
rect 20347 21732 20371 21734
rect 20427 21732 20451 21734
rect 20507 21732 20513 21734
rect 20205 21723 20513 21732
rect 19892 21004 19944 21010
rect 19892 20946 19944 20952
rect 20536 21004 20588 21010
rect 20536 20946 20588 20952
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18248 20602 18276 20742
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18340 20466 18368 20878
rect 18604 20868 18656 20874
rect 18604 20810 18656 20816
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18236 20324 18288 20330
rect 18236 20266 18288 20272
rect 18248 19854 18276 20266
rect 18340 19922 18368 20402
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18432 19990 18460 20334
rect 18420 19984 18472 19990
rect 18420 19926 18472 19932
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 17972 18414 18092 18442
rect 18156 18426 18184 18702
rect 18144 18420 18196 18426
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17420 16046 17448 18158
rect 17972 17338 18000 18414
rect 18144 18362 18196 18368
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18064 17882 18092 18226
rect 18432 18222 18460 19926
rect 18616 19854 18644 20810
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20602 18736 20742
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 19076 20330 19104 20810
rect 20205 20700 20513 20709
rect 20205 20698 20211 20700
rect 20267 20698 20291 20700
rect 20347 20698 20371 20700
rect 20427 20698 20451 20700
rect 20507 20698 20513 20700
rect 20267 20646 20269 20698
rect 20449 20646 20451 20698
rect 20205 20644 20211 20646
rect 20267 20644 20291 20646
rect 20347 20644 20371 20646
rect 20427 20644 20451 20646
rect 20507 20644 20513 20646
rect 20205 20635 20513 20644
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18892 19854 18920 20198
rect 19545 20156 19853 20165
rect 19545 20154 19551 20156
rect 19607 20154 19631 20156
rect 19687 20154 19711 20156
rect 19767 20154 19791 20156
rect 19847 20154 19853 20156
rect 19607 20102 19609 20154
rect 19789 20102 19791 20154
rect 19545 20100 19551 20102
rect 19607 20100 19631 20102
rect 19687 20100 19711 20102
rect 19767 20100 19791 20102
rect 19847 20100 19853 20102
rect 19545 20091 19853 20100
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18524 17678 18552 19654
rect 20205 19612 20513 19621
rect 20205 19610 20211 19612
rect 20267 19610 20291 19612
rect 20347 19610 20371 19612
rect 20427 19610 20451 19612
rect 20507 19610 20513 19612
rect 20267 19558 20269 19610
rect 20449 19558 20451 19610
rect 20205 19556 20211 19558
rect 20267 19556 20291 19558
rect 20347 19556 20371 19558
rect 20427 19556 20451 19558
rect 20507 19556 20513 19558
rect 20205 19547 20513 19556
rect 19545 19068 19853 19077
rect 19545 19066 19551 19068
rect 19607 19066 19631 19068
rect 19687 19066 19711 19068
rect 19767 19066 19791 19068
rect 19847 19066 19853 19068
rect 19607 19014 19609 19066
rect 19789 19014 19791 19066
rect 19545 19012 19551 19014
rect 19607 19012 19631 19014
rect 19687 19012 19711 19014
rect 19767 19012 19791 19014
rect 19847 19012 19853 19014
rect 19545 19003 19853 19012
rect 20205 18524 20513 18533
rect 20205 18522 20211 18524
rect 20267 18522 20291 18524
rect 20347 18522 20371 18524
rect 20427 18522 20451 18524
rect 20507 18522 20513 18524
rect 20267 18470 20269 18522
rect 20449 18470 20451 18522
rect 20205 18468 20211 18470
rect 20267 18468 20291 18470
rect 20347 18468 20371 18470
rect 20427 18468 20451 18470
rect 20507 18468 20513 18470
rect 20205 18459 20513 18468
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 18524 17134 18552 17614
rect 18616 17202 18644 17682
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 19064 17604 19116 17610
rect 19064 17546 19116 17552
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18708 16574 18736 17478
rect 18800 17338 18828 17546
rect 19076 17338 19104 17546
rect 19352 17338 19380 18294
rect 19444 17728 19472 18294
rect 19545 17980 19853 17989
rect 19545 17978 19551 17980
rect 19607 17978 19631 17980
rect 19687 17978 19711 17980
rect 19767 17978 19791 17980
rect 19847 17978 19853 17980
rect 19607 17926 19609 17978
rect 19789 17926 19791 17978
rect 19545 17924 19551 17926
rect 19607 17924 19631 17926
rect 19687 17924 19711 17926
rect 19767 17924 19791 17926
rect 19847 17924 19853 17926
rect 19545 17915 19853 17924
rect 19524 17740 19576 17746
rect 19444 17700 19524 17728
rect 19524 17682 19576 17688
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19536 17202 19564 17682
rect 19904 17678 19932 18294
rect 20548 18222 20576 20946
rect 22008 20936 22060 20942
rect 22008 20878 22060 20884
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21836 20466 21864 20742
rect 22020 20505 22048 20878
rect 22006 20496 22062 20505
rect 21824 20460 21876 20466
rect 22006 20431 22062 20440
rect 21824 20402 21876 20408
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19904 17134 19932 17614
rect 20205 17436 20513 17445
rect 20205 17434 20211 17436
rect 20267 17434 20291 17436
rect 20347 17434 20371 17436
rect 20427 17434 20451 17436
rect 20507 17434 20513 17436
rect 20267 17382 20269 17434
rect 20449 17382 20451 17434
rect 20205 17380 20211 17382
rect 20267 17380 20291 17382
rect 20347 17380 20371 17382
rect 20427 17380 20451 17382
rect 20507 17380 20513 17382
rect 20205 17371 20513 17380
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19545 16892 19853 16901
rect 19545 16890 19551 16892
rect 19607 16890 19631 16892
rect 19687 16890 19711 16892
rect 19767 16890 19791 16892
rect 19847 16890 19853 16892
rect 19607 16838 19609 16890
rect 19789 16838 19791 16890
rect 19545 16836 19551 16838
rect 19607 16836 19631 16838
rect 19687 16836 19711 16838
rect 19767 16836 19791 16838
rect 19847 16836 19853 16838
rect 19545 16827 19853 16836
rect 18708 16546 18828 16574
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 18340 15162 18368 16050
rect 18432 15706 18460 16050
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18800 15502 18828 16546
rect 20205 16348 20513 16357
rect 20205 16346 20211 16348
rect 20267 16346 20291 16348
rect 20347 16346 20371 16348
rect 20427 16346 20451 16348
rect 20507 16346 20513 16348
rect 20267 16294 20269 16346
rect 20449 16294 20451 16346
rect 20205 16292 20211 16294
rect 20267 16292 20291 16294
rect 20347 16292 20371 16294
rect 20427 16292 20451 16294
rect 20507 16292 20513 16294
rect 20205 16283 20513 16292
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18892 14958 18920 15914
rect 19545 15804 19853 15813
rect 19545 15802 19551 15804
rect 19607 15802 19631 15804
rect 19687 15802 19711 15804
rect 19767 15802 19791 15804
rect 19847 15802 19853 15804
rect 19607 15750 19609 15802
rect 19789 15750 19791 15802
rect 19545 15748 19551 15750
rect 19607 15748 19631 15750
rect 19687 15748 19711 15750
rect 19767 15748 19791 15750
rect 19847 15748 19853 15750
rect 19545 15739 19853 15748
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19168 14958 19196 15506
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19260 14618 19288 14962
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19352 14414 19380 15642
rect 20205 15260 20513 15269
rect 20205 15258 20211 15260
rect 20267 15258 20291 15260
rect 20347 15258 20371 15260
rect 20427 15258 20451 15260
rect 20507 15258 20513 15260
rect 20267 15206 20269 15258
rect 20449 15206 20451 15258
rect 20205 15204 20211 15206
rect 20267 15204 20291 15206
rect 20347 15204 20371 15206
rect 20427 15204 20451 15206
rect 20507 15204 20513 15206
rect 20205 15195 20513 15204
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 19444 14550 19472 15030
rect 20548 15026 20576 18158
rect 20640 17746 20668 20334
rect 22008 19848 22060 19854
rect 22006 19816 22008 19825
rect 22060 19816 22062 19825
rect 22006 19751 22062 19760
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 21008 18290 21036 18566
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 19892 14884 19944 14890
rect 19892 14826 19944 14832
rect 19545 14716 19853 14725
rect 19545 14714 19551 14716
rect 19607 14714 19631 14716
rect 19687 14714 19711 14716
rect 19767 14714 19791 14716
rect 19847 14714 19853 14716
rect 19607 14662 19609 14714
rect 19789 14662 19791 14714
rect 19545 14660 19551 14662
rect 19607 14660 19631 14662
rect 19687 14660 19711 14662
rect 19767 14660 19791 14662
rect 19847 14660 19853 14662
rect 19545 14651 19853 14660
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 17328 14278 17356 14350
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17328 14074 17356 14214
rect 18892 14074 18920 14282
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 19444 13870 19472 14486
rect 19904 14414 19932 14826
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 13938 19932 14350
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15856 11354 15884 11698
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15948 11150 15976 11698
rect 16960 11694 16988 12038
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16224 11218 16252 11494
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 16500 10810 16528 11222
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 16684 10062 16712 11494
rect 16960 10130 16988 11630
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16868 9654 16896 9862
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 9042 15608 9318
rect 16776 9042 16804 9522
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15304 7886 15332 8434
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 14832 7880 14884 7886
rect 14752 7828 14832 7834
rect 14752 7822 14884 7828
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 14752 7806 14872 7822
rect 14752 7410 14780 7806
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 14892 7644 15200 7653
rect 14892 7642 14898 7644
rect 14954 7642 14978 7644
rect 15034 7642 15058 7644
rect 15114 7642 15138 7644
rect 15194 7642 15200 7644
rect 14954 7590 14956 7642
rect 15136 7590 15138 7642
rect 14892 7588 14898 7590
rect 14954 7588 14978 7590
rect 15034 7588 15058 7590
rect 15114 7588 15138 7590
rect 15194 7588 15200 7590
rect 14892 7579 15200 7588
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 15200 7404 15252 7410
rect 15304 7392 15332 7686
rect 15252 7364 15332 7392
rect 15200 7346 15252 7352
rect 15212 7002 15240 7346
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14892 6556 15200 6565
rect 14892 6554 14898 6556
rect 14954 6554 14978 6556
rect 15034 6554 15058 6556
rect 15114 6554 15138 6556
rect 15194 6554 15200 6556
rect 14954 6502 14956 6554
rect 15136 6502 15138 6554
rect 14892 6500 14898 6502
rect 14954 6500 14978 6502
rect 15034 6500 15058 6502
rect 15114 6500 15138 6502
rect 15194 6500 15200 6502
rect 14892 6491 15200 6500
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14232 6012 14540 6021
rect 14232 6010 14238 6012
rect 14294 6010 14318 6012
rect 14374 6010 14398 6012
rect 14454 6010 14478 6012
rect 14534 6010 14540 6012
rect 14294 5958 14296 6010
rect 14476 5958 14478 6010
rect 14232 5956 14238 5958
rect 14294 5956 14318 5958
rect 14374 5956 14398 5958
rect 14454 5956 14478 5958
rect 14534 5956 14540 5958
rect 14232 5947 14540 5956
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13832 4678 13952 4706
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 13556 4282 13584 4490
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13556 3466 13584 4082
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13648 3534 13676 4014
rect 13832 3738 13860 4218
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13556 3194 13584 3402
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13832 2582 13860 2994
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13924 2446 13952 4678
rect 14016 4146 14044 5782
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14004 4004 14056 4010
rect 14004 3946 14056 3952
rect 14016 3738 14044 3946
rect 14108 3942 14136 5170
rect 14232 4924 14540 4933
rect 14232 4922 14238 4924
rect 14294 4922 14318 4924
rect 14374 4922 14398 4924
rect 14454 4922 14478 4924
rect 14534 4922 14540 4924
rect 14294 4870 14296 4922
rect 14476 4870 14478 4922
rect 14232 4868 14238 4870
rect 14294 4868 14318 4870
rect 14374 4868 14398 4870
rect 14454 4868 14478 4870
rect 14534 4868 14540 4870
rect 14232 4859 14540 4868
rect 14568 4010 14596 6190
rect 14660 5914 14688 6326
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14936 5778 14964 6054
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14660 4690 14688 5102
rect 14752 4826 14780 5510
rect 14892 5468 15200 5477
rect 14892 5466 14898 5468
rect 14954 5466 14978 5468
rect 15034 5466 15058 5468
rect 15114 5466 15138 5468
rect 15194 5466 15200 5468
rect 14954 5414 14956 5466
rect 15136 5414 15138 5466
rect 14892 5412 14898 5414
rect 14954 5412 14978 5414
rect 15034 5412 15058 5414
rect 15114 5412 15138 5414
rect 15194 5412 15200 5414
rect 14892 5403 15200 5412
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 15120 4554 15148 5170
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 14892 4380 15200 4389
rect 14892 4378 14898 4380
rect 14954 4378 14978 4380
rect 15034 4378 15058 4380
rect 15114 4378 15138 4380
rect 15194 4378 15200 4380
rect 14954 4326 14956 4378
rect 15136 4326 15138 4378
rect 14892 4324 14898 4326
rect 14954 4324 14978 4326
rect 15034 4324 15058 4326
rect 15114 4324 15138 4326
rect 15194 4324 15200 4326
rect 14892 4315 15200 4324
rect 15488 4146 15516 4422
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14232 3836 14540 3845
rect 14232 3834 14238 3836
rect 14294 3834 14318 3836
rect 14374 3834 14398 3836
rect 14454 3834 14478 3836
rect 14534 3834 14540 3836
rect 14294 3782 14296 3834
rect 14476 3782 14478 3834
rect 14232 3780 14238 3782
rect 14294 3780 14318 3782
rect 14374 3780 14398 3782
rect 14454 3780 14478 3782
rect 14534 3780 14540 3782
rect 14232 3771 14540 3780
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14200 3058 14228 3470
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 3194 14320 3334
rect 14660 3194 14688 3402
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14892 3292 15200 3301
rect 14892 3290 14898 3292
rect 14954 3290 14978 3292
rect 15034 3290 15058 3292
rect 15114 3290 15138 3292
rect 15194 3290 15200 3292
rect 14954 3238 14956 3290
rect 15136 3238 15138 3290
rect 14892 3236 14898 3238
rect 14954 3236 14978 3238
rect 15034 3236 15058 3238
rect 15114 3236 15138 3238
rect 15194 3236 15200 3238
rect 14892 3227 15200 3236
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 14200 2854 14228 2994
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14232 2748 14540 2757
rect 14232 2746 14238 2748
rect 14294 2746 14318 2748
rect 14374 2746 14398 2748
rect 14454 2746 14478 2748
rect 14534 2746 14540 2748
rect 14294 2694 14296 2746
rect 14476 2694 14478 2746
rect 14232 2692 14238 2694
rect 14294 2692 14318 2694
rect 14374 2692 14398 2694
rect 14454 2692 14478 2694
rect 14534 2692 14540 2694
rect 14232 2683 14540 2692
rect 14936 2650 14964 2790
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15028 2582 15056 2994
rect 15304 2990 15332 3334
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 15580 2446 15608 7142
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15856 4622 15884 6802
rect 16132 6390 16160 6802
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16132 3602 16160 4082
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16224 2446 16252 8298
rect 16960 7954 16988 10066
rect 17144 9738 17172 13738
rect 19545 13628 19853 13637
rect 19545 13626 19551 13628
rect 19607 13626 19631 13628
rect 19687 13626 19711 13628
rect 19767 13626 19791 13628
rect 19847 13626 19853 13628
rect 19607 13574 19609 13626
rect 19789 13574 19791 13626
rect 19545 13572 19551 13574
rect 19607 13572 19631 13574
rect 19687 13572 19711 13574
rect 19767 13572 19791 13574
rect 19847 13572 19853 13574
rect 19545 13563 19853 13572
rect 20088 13394 20116 14962
rect 20640 14958 20668 17682
rect 21100 16590 21128 18226
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21560 17785 21588 18022
rect 21546 17776 21602 17785
rect 21546 17711 21602 17720
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21376 16522 21404 17138
rect 21546 17096 21602 17105
rect 21546 17031 21548 17040
rect 21600 17031 21602 17040
rect 21548 17002 21600 17008
rect 21364 16516 21416 16522
rect 21364 16458 21416 16464
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15502 21128 15846
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21100 15162 21128 15438
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21192 15162 21220 15302
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20364 14618 20392 14894
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20205 14172 20513 14181
rect 20205 14170 20211 14172
rect 20267 14170 20291 14172
rect 20347 14170 20371 14172
rect 20427 14170 20451 14172
rect 20507 14170 20513 14172
rect 20267 14118 20269 14170
rect 20449 14118 20451 14170
rect 20205 14116 20211 14118
rect 20267 14116 20291 14118
rect 20347 14116 20371 14118
rect 20427 14116 20451 14118
rect 20507 14116 20513 14118
rect 20205 14107 20513 14116
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19628 12918 19656 13126
rect 20205 13084 20513 13093
rect 20205 13082 20211 13084
rect 20267 13082 20291 13084
rect 20347 13082 20371 13084
rect 20427 13082 20451 13084
rect 20507 13082 20513 13084
rect 20267 13030 20269 13082
rect 20449 13030 20451 13082
rect 20205 13028 20211 13030
rect 20267 13028 20291 13030
rect 20347 13028 20371 13030
rect 20427 13028 20451 13030
rect 20507 13028 20513 13030
rect 20205 13019 20513 13028
rect 20548 12918 20576 14214
rect 20640 13802 20668 14894
rect 20732 14414 20760 15030
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 21652 14006 21680 19450
rect 21836 17678 21864 19654
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22020 19145 22048 19314
rect 22006 19136 22062 19145
rect 22006 19071 22062 19080
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22020 18465 22048 18702
rect 22006 18456 22062 18465
rect 22006 18391 22062 18400
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 21732 16448 21784 16454
rect 22020 16425 22048 16526
rect 21732 16390 21784 16396
rect 22006 16416 22062 16425
rect 21640 14000 21692 14006
rect 21640 13942 21692 13948
rect 20628 13796 20680 13802
rect 20628 13738 20680 13744
rect 21744 13326 21772 16390
rect 22006 16351 22062 16360
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22020 15745 22048 16050
rect 22006 15736 22062 15745
rect 22006 15671 22062 15680
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21824 15360 21876 15366
rect 21824 15302 21876 15308
rect 21836 15094 21864 15302
rect 21824 15088 21876 15094
rect 22020 15065 22048 15438
rect 21824 15030 21876 15036
rect 22006 15056 22062 15065
rect 22006 14991 22062 15000
rect 22008 14408 22060 14414
rect 22006 14376 22008 14385
rect 22060 14376 22062 14385
rect 22006 14311 22062 14320
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21824 13728 21876 13734
rect 22020 13705 22048 13874
rect 21824 13670 21876 13676
rect 22006 13696 22062 13705
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21836 12986 21864 13670
rect 22006 13631 22062 13640
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22020 13025 22048 13262
rect 22006 13016 22062 13025
rect 21824 12980 21876 12986
rect 22006 12951 22062 12960
rect 21824 12922 21876 12928
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19616 12912 19668 12918
rect 20536 12912 20588 12918
rect 19616 12854 19668 12860
rect 20456 12860 20536 12866
rect 20456 12854 20588 12860
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17696 11218 17724 12242
rect 18064 12238 18092 12650
rect 18248 12306 18276 12718
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17880 11898 17908 12106
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18064 11830 18092 12038
rect 18248 11830 18276 12242
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11898 18368 12038
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18156 11354 18184 11698
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 18432 11064 18460 12582
rect 18524 12238 18552 12582
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18616 11830 18644 12650
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18708 11694 18736 12242
rect 19352 12238 19380 12854
rect 20456 12838 20576 12854
rect 22008 12844 22060 12850
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19444 12442 19472 12718
rect 19545 12540 19853 12549
rect 19545 12538 19551 12540
rect 19607 12538 19631 12540
rect 19687 12538 19711 12540
rect 19767 12538 19791 12540
rect 19847 12538 19853 12540
rect 19607 12486 19609 12538
rect 19789 12486 19791 12538
rect 19545 12484 19551 12486
rect 19607 12484 19631 12486
rect 19687 12484 19711 12486
rect 19767 12484 19791 12486
rect 19847 12484 19853 12486
rect 19545 12475 19853 12484
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19904 12306 19932 12718
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 20456 12238 20484 12838
rect 22008 12786 22060 12792
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20548 12442 20576 12718
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20205 11996 20513 12005
rect 20205 11994 20211 11996
rect 20267 11994 20291 11996
rect 20347 11994 20371 11996
rect 20427 11994 20451 11996
rect 20507 11994 20513 11996
rect 20267 11942 20269 11994
rect 20449 11942 20451 11994
rect 20205 11940 20211 11942
rect 20267 11940 20291 11942
rect 20347 11940 20371 11942
rect 20427 11940 20451 11942
rect 20507 11940 20513 11942
rect 20205 11931 20513 11940
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18512 11076 18564 11082
rect 18432 11036 18512 11064
rect 18512 11018 18564 11024
rect 18708 10266 18736 11630
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 19545 11452 19853 11461
rect 19545 11450 19551 11452
rect 19607 11450 19631 11452
rect 19687 11450 19711 11452
rect 19767 11450 19791 11452
rect 19847 11450 19853 11452
rect 19607 11398 19609 11450
rect 19789 11398 19791 11450
rect 19545 11396 19551 11398
rect 19607 11396 19631 11398
rect 19687 11396 19711 11398
rect 19767 11396 19791 11398
rect 19847 11396 19853 11398
rect 19545 11387 19853 11396
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17052 9710 17172 9738
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16408 3534 16436 4014
rect 16592 3942 16620 6666
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 6458 16712 6598
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16684 4622 16712 5102
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16684 4078 16712 4558
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16500 3194 16528 3538
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16776 2446 16804 7210
rect 16960 6866 16988 7890
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17052 6474 17080 9710
rect 17880 9586 17908 9998
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17144 8498 17172 9522
rect 18064 9518 18092 9862
rect 18156 9586 18184 9862
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18432 9110 18460 10066
rect 18708 10062 18736 10202
rect 19076 10130 19104 10950
rect 20205 10908 20513 10917
rect 20205 10906 20211 10908
rect 20267 10906 20291 10908
rect 20347 10906 20371 10908
rect 20427 10906 20451 10908
rect 20507 10906 20513 10908
rect 20267 10854 20269 10906
rect 20449 10854 20451 10906
rect 20205 10852 20211 10854
rect 20267 10852 20291 10854
rect 20347 10852 20371 10854
rect 20427 10852 20451 10854
rect 20507 10852 20513 10854
rect 20205 10843 20513 10852
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 18892 9586 18920 9862
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 19352 9518 19380 10610
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19444 10130 19472 10406
rect 19545 10364 19853 10373
rect 19545 10362 19551 10364
rect 19607 10362 19631 10364
rect 19687 10362 19711 10364
rect 19767 10362 19791 10364
rect 19847 10362 19853 10364
rect 19607 10310 19609 10362
rect 19789 10310 19791 10362
rect 19545 10308 19551 10310
rect 19607 10308 19631 10310
rect 19687 10308 19711 10310
rect 19767 10308 19791 10310
rect 19847 10308 19853 10310
rect 19545 10299 19853 10308
rect 19996 10266 20024 10474
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19536 9586 19564 10202
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19628 9722 19656 9862
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 20088 9602 20116 10406
rect 20456 10062 20484 10610
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20548 10130 20576 10406
rect 20640 10130 20668 11494
rect 20732 10810 20760 12718
rect 22020 12345 22048 12786
rect 22006 12336 22062 12345
rect 22006 12271 22062 12280
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22020 11665 22048 11698
rect 22006 11656 22062 11665
rect 22006 11591 22062 11600
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22020 10985 22048 11086
rect 22006 10976 22062 10985
rect 22006 10911 22062 10920
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20732 10130 20760 10746
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22020 10305 22048 10610
rect 22006 10296 22062 10305
rect 22006 10231 22062 10240
rect 21180 10192 21232 10198
rect 21180 10134 21232 10140
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20444 10056 20496 10062
rect 20640 10010 20668 10066
rect 20444 9998 20496 10004
rect 20548 9982 20668 10010
rect 20205 9820 20513 9829
rect 20205 9818 20211 9820
rect 20267 9818 20291 9820
rect 20347 9818 20371 9820
rect 20427 9818 20451 9820
rect 20507 9818 20513 9820
rect 20267 9766 20269 9818
rect 20449 9766 20451 9818
rect 20205 9764 20211 9766
rect 20267 9764 20291 9766
rect 20347 9764 20371 9766
rect 20427 9764 20451 9766
rect 20507 9764 20513 9766
rect 20205 9755 20513 9764
rect 20168 9648 20220 9654
rect 20088 9596 20168 9602
rect 20088 9590 20220 9596
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19892 9580 19944 9586
rect 20088 9574 20208 9590
rect 19892 9522 19944 9528
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18800 9042 18828 9454
rect 19545 9276 19853 9285
rect 19545 9274 19551 9276
rect 19607 9274 19631 9276
rect 19687 9274 19711 9276
rect 19767 9274 19791 9276
rect 19847 9274 19853 9276
rect 19607 9222 19609 9274
rect 19789 9222 19791 9274
rect 19545 9220 19551 9222
rect 19607 9220 19631 9222
rect 19687 9220 19711 9222
rect 19767 9220 19791 9222
rect 19847 9220 19853 9222
rect 19545 9211 19853 9220
rect 19904 9178 19932 9522
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 19996 8498 20024 9318
rect 20205 8732 20513 8741
rect 20205 8730 20211 8732
rect 20267 8730 20291 8732
rect 20347 8730 20371 8732
rect 20427 8730 20451 8732
rect 20507 8730 20513 8732
rect 20267 8678 20269 8730
rect 20449 8678 20451 8730
rect 20205 8676 20211 8678
rect 20267 8676 20291 8678
rect 20347 8676 20371 8678
rect 20427 8676 20451 8678
rect 20507 8676 20513 8678
rect 20205 8667 20513 8676
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 17144 6662 17172 8434
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 17604 7954 17632 8230
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17868 7880 17920 7886
rect 17920 7828 18184 7834
rect 17868 7822 18184 7828
rect 17236 6934 17264 7822
rect 17880 7818 18184 7822
rect 17880 7812 18196 7818
rect 17880 7806 18144 7812
rect 18144 7754 18196 7760
rect 18984 7478 19012 8230
rect 19260 7954 19288 8366
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 19260 7342 19288 7890
rect 19444 7886 19472 8230
rect 19545 8188 19853 8197
rect 19545 8186 19551 8188
rect 19607 8186 19631 8188
rect 19687 8186 19711 8188
rect 19767 8186 19791 8188
rect 19847 8186 19853 8188
rect 19607 8134 19609 8186
rect 19789 8134 19791 8186
rect 19545 8132 19551 8134
rect 19607 8132 19631 8134
rect 19687 8132 19711 8134
rect 19767 8132 19791 8134
rect 19847 8132 19853 8134
rect 19545 8123 19853 8132
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19628 7546 19656 7686
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17052 6446 17172 6474
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17052 5166 17080 6258
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 16960 3738 16988 4490
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17052 3738 17080 4082
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16856 3528 16908 3534
rect 17144 3482 17172 6446
rect 17236 6254 17264 6870
rect 18340 6866 18368 7142
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17236 5302 17264 6190
rect 18248 5370 18276 6666
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18432 6254 18460 6598
rect 18800 6322 18828 6598
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17236 4214 17264 5238
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17696 4826 17724 5170
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17880 4826 17908 5102
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 18708 4622 18736 5510
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 16856 3470 16908 3476
rect 16868 3194 16896 3470
rect 17052 3466 17172 3482
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17040 3460 17172 3466
rect 17092 3454 17172 3460
rect 17040 3402 17092 3408
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17328 3058 17356 3470
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17880 3194 17908 3334
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17052 2650 17080 2994
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 18800 2446 18828 6122
rect 18892 5710 18920 6190
rect 19076 5846 19104 6802
rect 19352 6458 19380 7414
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19444 6798 19472 7210
rect 19545 7100 19853 7109
rect 19545 7098 19551 7100
rect 19607 7098 19631 7100
rect 19687 7098 19711 7100
rect 19767 7098 19791 7100
rect 19847 7098 19853 7100
rect 19607 7046 19609 7098
rect 19789 7046 19791 7098
rect 19545 7044 19551 7046
rect 19607 7044 19631 7046
rect 19687 7044 19711 7046
rect 19767 7044 19791 7046
rect 19847 7044 19853 7046
rect 19545 7035 19853 7044
rect 19904 7002 19932 7686
rect 20205 7644 20513 7653
rect 20205 7642 20211 7644
rect 20267 7642 20291 7644
rect 20347 7642 20371 7644
rect 20427 7642 20451 7644
rect 20507 7642 20513 7644
rect 20267 7590 20269 7642
rect 20449 7590 20451 7642
rect 20205 7588 20211 7590
rect 20267 7588 20291 7590
rect 20347 7588 20371 7590
rect 20427 7588 20451 7590
rect 20507 7588 20513 7590
rect 20205 7579 20513 7588
rect 20548 7342 20576 9982
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20640 9518 20668 9862
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19545 6012 19853 6021
rect 19545 6010 19551 6012
rect 19607 6010 19631 6012
rect 19687 6010 19711 6012
rect 19767 6010 19791 6012
rect 19847 6010 19853 6012
rect 19607 5958 19609 6010
rect 19789 5958 19791 6010
rect 19545 5956 19551 5958
rect 19607 5956 19631 5958
rect 19687 5956 19711 5958
rect 19767 5956 19791 5958
rect 19847 5956 19853 5958
rect 19545 5947 19853 5956
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18892 5166 18920 5646
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 19168 4758 19196 5170
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19260 4826 19288 5034
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 19168 4622 19196 4694
rect 19352 4690 19380 5102
rect 19545 4924 19853 4933
rect 19545 4922 19551 4924
rect 19607 4922 19631 4924
rect 19687 4922 19711 4924
rect 19767 4922 19791 4924
rect 19847 4922 19853 4924
rect 19607 4870 19609 4922
rect 19789 4870 19791 4922
rect 19545 4868 19551 4870
rect 19607 4868 19631 4870
rect 19687 4868 19711 4870
rect 19767 4868 19791 4870
rect 19847 4868 19853 4870
rect 19545 4859 19853 4868
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19168 4298 19196 4558
rect 19352 4554 19380 4626
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19076 4282 19196 4298
rect 19064 4276 19196 4282
rect 19116 4270 19196 4276
rect 19064 4218 19116 4224
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19260 3738 19288 4014
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19352 3126 19380 4014
rect 19444 3534 19472 4150
rect 19996 4078 20024 7278
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20272 6798 20300 7210
rect 20732 6934 20760 10066
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20720 6928 20772 6934
rect 20720 6870 20772 6876
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20088 6322 20116 6734
rect 20205 6556 20513 6565
rect 20205 6554 20211 6556
rect 20267 6554 20291 6556
rect 20347 6554 20371 6556
rect 20427 6554 20451 6556
rect 20507 6554 20513 6556
rect 20267 6502 20269 6554
rect 20449 6502 20451 6554
rect 20205 6500 20211 6502
rect 20267 6500 20291 6502
rect 20347 6500 20371 6502
rect 20427 6500 20451 6502
rect 20507 6500 20513 6502
rect 20205 6491 20513 6500
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 20548 6254 20576 6734
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20205 5468 20513 5477
rect 20205 5466 20211 5468
rect 20267 5466 20291 5468
rect 20347 5466 20371 5468
rect 20427 5466 20451 5468
rect 20507 5466 20513 5468
rect 20267 5414 20269 5466
rect 20449 5414 20451 5466
rect 20205 5412 20211 5414
rect 20267 5412 20291 5414
rect 20347 5412 20371 5414
rect 20427 5412 20451 5414
rect 20507 5412 20513 5414
rect 20205 5403 20513 5412
rect 20732 4690 20760 6870
rect 20916 6866 20944 7142
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21192 6322 21220 10134
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21284 9586 21312 9862
rect 21376 9722 21404 9862
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21744 9654 21772 9998
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21732 9648 21784 9654
rect 21928 9625 21956 9862
rect 21732 9590 21784 9596
rect 21914 9616 21970 9625
rect 21272 9580 21324 9586
rect 21914 9551 21970 9560
rect 21272 9522 21324 9528
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21284 5370 21312 9522
rect 21914 8936 21970 8945
rect 21914 8871 21970 8880
rect 21928 8838 21956 8871
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21548 8356 21600 8362
rect 21548 8298 21600 8304
rect 21560 8265 21588 8298
rect 21546 8256 21602 8265
rect 21546 8191 21602 8200
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21928 7585 21956 7686
rect 21914 7576 21970 7585
rect 21914 7511 21970 7520
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 21836 6662 21864 7346
rect 22020 6905 22048 7346
rect 22006 6896 22062 6905
rect 22006 6831 22062 6840
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21546 6216 21602 6225
rect 21546 6151 21548 6160
rect 21600 6151 21602 6160
rect 21548 6122 21600 6128
rect 21836 5914 21864 6598
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 22008 5704 22060 5710
rect 22008 5646 22060 5652
rect 22020 5545 22048 5646
rect 22006 5536 22062 5545
rect 22006 5471 22062 5480
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 22020 4865 22048 5170
rect 22006 4856 22062 4865
rect 22006 4791 22062 4800
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20205 4380 20513 4389
rect 20205 4378 20211 4380
rect 20267 4378 20291 4380
rect 20347 4378 20371 4380
rect 20427 4378 20451 4380
rect 20507 4378 20513 4380
rect 20267 4326 20269 4378
rect 20449 4326 20451 4378
rect 20205 4324 20211 4326
rect 20267 4324 20291 4326
rect 20347 4324 20371 4326
rect 20427 4324 20451 4326
rect 20507 4324 20513 4326
rect 20205 4315 20513 4324
rect 20732 4162 20760 4626
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22020 4185 22048 4558
rect 20640 4134 20760 4162
rect 22006 4176 22062 4185
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19545 3836 19853 3845
rect 19545 3834 19551 3836
rect 19607 3834 19631 3836
rect 19687 3834 19711 3836
rect 19767 3834 19791 3836
rect 19847 3834 19853 3836
rect 19607 3782 19609 3834
rect 19789 3782 19791 3834
rect 19545 3780 19551 3782
rect 19607 3780 19631 3782
rect 19687 3780 19711 3782
rect 19767 3780 19791 3782
rect 19847 3780 19853 3782
rect 19545 3771 19853 3780
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19444 2650 19472 3470
rect 20205 3292 20513 3301
rect 20205 3290 20211 3292
rect 20267 3290 20291 3292
rect 20347 3290 20371 3292
rect 20427 3290 20451 3292
rect 20507 3290 20513 3292
rect 20267 3238 20269 3290
rect 20449 3238 20451 3290
rect 20205 3236 20211 3238
rect 20267 3236 20291 3238
rect 20347 3236 20371 3238
rect 20427 3236 20451 3238
rect 20507 3236 20513 3238
rect 20205 3227 20513 3236
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19545 2748 19853 2757
rect 19545 2746 19551 2748
rect 19607 2746 19631 2748
rect 19687 2746 19711 2748
rect 19767 2746 19791 2748
rect 19847 2746 19853 2748
rect 19607 2694 19609 2746
rect 19789 2694 19791 2746
rect 19545 2692 19551 2694
rect 19607 2692 19631 2694
rect 19687 2692 19711 2694
rect 19767 2692 19791 2694
rect 19847 2692 19853 2694
rect 19545 2683 19853 2692
rect 20088 2650 20116 2994
rect 20640 2990 20668 4134
rect 22006 4111 22062 4120
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 12268 800 12296 2382
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 12912 800 12940 2314
rect 13556 800 13584 2382
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 800 14228 2246
rect 14752 1306 14780 2382
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 14892 2204 15200 2213
rect 14892 2202 14898 2204
rect 14954 2202 14978 2204
rect 15034 2202 15058 2204
rect 15114 2202 15138 2204
rect 15194 2202 15200 2204
rect 14954 2150 14956 2202
rect 15136 2150 15138 2202
rect 14892 2148 14898 2150
rect 14954 2148 14978 2150
rect 15034 2148 15058 2150
rect 15114 2148 15138 2150
rect 15194 2148 15200 2150
rect 14892 2139 15200 2148
rect 14752 1278 14872 1306
rect 14844 800 14872 1278
rect 15488 800 15516 2246
rect 16132 800 16160 2246
rect 16776 800 16804 2246
rect 17420 800 17448 2382
rect 18064 800 18092 2382
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18708 800 18736 2246
rect 19352 800 19380 2382
rect 19996 800 20024 2382
rect 20205 2204 20513 2213
rect 20205 2202 20211 2204
rect 20267 2202 20291 2204
rect 20347 2202 20371 2204
rect 20427 2202 20451 2204
rect 20507 2202 20513 2204
rect 20267 2150 20269 2202
rect 20449 2150 20451 2202
rect 20205 2148 20211 2150
rect 20267 2148 20291 2150
rect 20347 2148 20371 2150
rect 20427 2148 20451 2150
rect 20507 2148 20513 2150
rect 20205 2139 20513 2148
rect 9784 734 9996 762
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
<< via2 >>
rect 3612 23418 3668 23420
rect 3692 23418 3748 23420
rect 3772 23418 3828 23420
rect 3852 23418 3908 23420
rect 3612 23366 3658 23418
rect 3658 23366 3668 23418
rect 3692 23366 3722 23418
rect 3722 23366 3734 23418
rect 3734 23366 3748 23418
rect 3772 23366 3786 23418
rect 3786 23366 3798 23418
rect 3798 23366 3828 23418
rect 3852 23366 3862 23418
rect 3862 23366 3908 23418
rect 3612 23364 3668 23366
rect 3692 23364 3748 23366
rect 3772 23364 3828 23366
rect 3852 23364 3908 23366
rect 8925 23418 8981 23420
rect 9005 23418 9061 23420
rect 9085 23418 9141 23420
rect 9165 23418 9221 23420
rect 8925 23366 8971 23418
rect 8971 23366 8981 23418
rect 9005 23366 9035 23418
rect 9035 23366 9047 23418
rect 9047 23366 9061 23418
rect 9085 23366 9099 23418
rect 9099 23366 9111 23418
rect 9111 23366 9141 23418
rect 9165 23366 9175 23418
rect 9175 23366 9221 23418
rect 8925 23364 8981 23366
rect 9005 23364 9061 23366
rect 9085 23364 9141 23366
rect 9165 23364 9221 23366
rect 4272 22874 4328 22876
rect 4352 22874 4408 22876
rect 4432 22874 4488 22876
rect 4512 22874 4568 22876
rect 4272 22822 4318 22874
rect 4318 22822 4328 22874
rect 4352 22822 4382 22874
rect 4382 22822 4394 22874
rect 4394 22822 4408 22874
rect 4432 22822 4446 22874
rect 4446 22822 4458 22874
rect 4458 22822 4488 22874
rect 4512 22822 4522 22874
rect 4522 22822 4568 22874
rect 4272 22820 4328 22822
rect 4352 22820 4408 22822
rect 4432 22820 4488 22822
rect 4512 22820 4568 22822
rect 846 22636 902 22672
rect 846 22616 848 22636
rect 848 22616 900 22636
rect 900 22616 902 22636
rect 846 21972 848 21992
rect 848 21972 900 21992
rect 900 21972 902 21992
rect 846 21936 902 21972
rect 846 21256 902 21312
rect 1490 20440 1546 20496
rect 846 19660 848 19680
rect 848 19660 900 19680
rect 900 19660 902 19680
rect 846 19624 902 19660
rect 1490 19116 1492 19136
rect 1492 19116 1544 19136
rect 1544 19116 1546 19136
rect 1490 19080 1546 19116
rect 846 18536 902 18592
rect 3612 22330 3668 22332
rect 3692 22330 3748 22332
rect 3772 22330 3828 22332
rect 3852 22330 3908 22332
rect 3612 22278 3658 22330
rect 3658 22278 3668 22330
rect 3692 22278 3722 22330
rect 3722 22278 3734 22330
rect 3734 22278 3748 22330
rect 3772 22278 3786 22330
rect 3786 22278 3798 22330
rect 3798 22278 3828 22330
rect 3852 22278 3862 22330
rect 3862 22278 3908 22330
rect 3612 22276 3668 22278
rect 3692 22276 3748 22278
rect 3772 22276 3828 22278
rect 3852 22276 3908 22278
rect 4272 21786 4328 21788
rect 4352 21786 4408 21788
rect 4432 21786 4488 21788
rect 4512 21786 4568 21788
rect 4272 21734 4318 21786
rect 4318 21734 4328 21786
rect 4352 21734 4382 21786
rect 4382 21734 4394 21786
rect 4394 21734 4408 21786
rect 4432 21734 4446 21786
rect 4446 21734 4458 21786
rect 4458 21734 4488 21786
rect 4512 21734 4522 21786
rect 4522 21734 4568 21786
rect 4272 21732 4328 21734
rect 4352 21732 4408 21734
rect 4432 21732 4488 21734
rect 4512 21732 4568 21734
rect 3612 21242 3668 21244
rect 3692 21242 3748 21244
rect 3772 21242 3828 21244
rect 3852 21242 3908 21244
rect 3612 21190 3658 21242
rect 3658 21190 3668 21242
rect 3692 21190 3722 21242
rect 3722 21190 3734 21242
rect 3734 21190 3748 21242
rect 3772 21190 3786 21242
rect 3786 21190 3798 21242
rect 3798 21190 3828 21242
rect 3852 21190 3862 21242
rect 3862 21190 3908 21242
rect 3612 21188 3668 21190
rect 3692 21188 3748 21190
rect 3772 21188 3828 21190
rect 3852 21188 3908 21190
rect 1490 17720 1546 17776
rect 846 16904 902 16960
rect 846 16532 848 16552
rect 848 16532 900 16552
rect 900 16532 902 16552
rect 846 16496 902 16532
rect 846 15852 848 15872
rect 848 15852 900 15872
rect 900 15852 902 15872
rect 846 15816 902 15852
rect 1398 15000 1454 15056
rect 846 14456 902 14512
rect 1398 13640 1454 13696
rect 846 13096 902 13152
rect 1398 12280 1454 12336
rect 846 11756 902 11792
rect 846 11736 848 11756
rect 848 11736 900 11756
rect 900 11736 902 11756
rect 1674 10920 1730 10976
rect 1490 10240 1546 10296
rect 1490 9560 1546 9616
rect 846 9052 848 9072
rect 848 9052 900 9072
rect 900 9052 902 9072
rect 846 9016 902 9052
rect 1490 8200 1546 8256
rect 3612 20154 3668 20156
rect 3692 20154 3748 20156
rect 3772 20154 3828 20156
rect 3852 20154 3908 20156
rect 3612 20102 3658 20154
rect 3658 20102 3668 20154
rect 3692 20102 3722 20154
rect 3722 20102 3734 20154
rect 3734 20102 3748 20154
rect 3772 20102 3786 20154
rect 3786 20102 3798 20154
rect 3798 20102 3828 20154
rect 3852 20102 3862 20154
rect 3862 20102 3908 20154
rect 3612 20100 3668 20102
rect 3692 20100 3748 20102
rect 3772 20100 3828 20102
rect 3852 20100 3908 20102
rect 4272 20698 4328 20700
rect 4352 20698 4408 20700
rect 4432 20698 4488 20700
rect 4512 20698 4568 20700
rect 4272 20646 4318 20698
rect 4318 20646 4328 20698
rect 4352 20646 4382 20698
rect 4382 20646 4394 20698
rect 4394 20646 4408 20698
rect 4432 20646 4446 20698
rect 4446 20646 4458 20698
rect 4458 20646 4488 20698
rect 4512 20646 4522 20698
rect 4522 20646 4568 20698
rect 4272 20644 4328 20646
rect 4352 20644 4408 20646
rect 4432 20644 4488 20646
rect 4512 20644 4568 20646
rect 4272 19610 4328 19612
rect 4352 19610 4408 19612
rect 4432 19610 4488 19612
rect 4512 19610 4568 19612
rect 4272 19558 4318 19610
rect 4318 19558 4328 19610
rect 4352 19558 4382 19610
rect 4382 19558 4394 19610
rect 4394 19558 4408 19610
rect 4432 19558 4446 19610
rect 4446 19558 4458 19610
rect 4458 19558 4488 19610
rect 4512 19558 4522 19610
rect 4522 19558 4568 19610
rect 4272 19556 4328 19558
rect 4352 19556 4408 19558
rect 4432 19556 4488 19558
rect 4512 19556 4568 19558
rect 3612 19066 3668 19068
rect 3692 19066 3748 19068
rect 3772 19066 3828 19068
rect 3852 19066 3908 19068
rect 3612 19014 3658 19066
rect 3658 19014 3668 19066
rect 3692 19014 3722 19066
rect 3722 19014 3734 19066
rect 3734 19014 3748 19066
rect 3772 19014 3786 19066
rect 3786 19014 3798 19066
rect 3798 19014 3828 19066
rect 3852 19014 3862 19066
rect 3862 19014 3908 19066
rect 3612 19012 3668 19014
rect 3692 19012 3748 19014
rect 3772 19012 3828 19014
rect 3852 19012 3908 19014
rect 4272 18522 4328 18524
rect 4352 18522 4408 18524
rect 4432 18522 4488 18524
rect 4512 18522 4568 18524
rect 4272 18470 4318 18522
rect 4318 18470 4328 18522
rect 4352 18470 4382 18522
rect 4382 18470 4394 18522
rect 4394 18470 4408 18522
rect 4432 18470 4446 18522
rect 4446 18470 4458 18522
rect 4458 18470 4488 18522
rect 4512 18470 4522 18522
rect 4522 18470 4568 18522
rect 4272 18468 4328 18470
rect 4352 18468 4408 18470
rect 4432 18468 4488 18470
rect 4512 18468 4568 18470
rect 3612 17978 3668 17980
rect 3692 17978 3748 17980
rect 3772 17978 3828 17980
rect 3852 17978 3908 17980
rect 3612 17926 3658 17978
rect 3658 17926 3668 17978
rect 3692 17926 3722 17978
rect 3722 17926 3734 17978
rect 3734 17926 3748 17978
rect 3772 17926 3786 17978
rect 3786 17926 3798 17978
rect 3798 17926 3828 17978
rect 3852 17926 3862 17978
rect 3862 17926 3908 17978
rect 3612 17924 3668 17926
rect 3692 17924 3748 17926
rect 3772 17924 3828 17926
rect 3852 17924 3908 17926
rect 3612 16890 3668 16892
rect 3692 16890 3748 16892
rect 3772 16890 3828 16892
rect 3852 16890 3908 16892
rect 3612 16838 3658 16890
rect 3658 16838 3668 16890
rect 3692 16838 3722 16890
rect 3722 16838 3734 16890
rect 3734 16838 3748 16890
rect 3772 16838 3786 16890
rect 3786 16838 3798 16890
rect 3798 16838 3828 16890
rect 3852 16838 3862 16890
rect 3862 16838 3908 16890
rect 3612 16836 3668 16838
rect 3692 16836 3748 16838
rect 3772 16836 3828 16838
rect 3852 16836 3908 16838
rect 4272 17434 4328 17436
rect 4352 17434 4408 17436
rect 4432 17434 4488 17436
rect 4512 17434 4568 17436
rect 4272 17382 4318 17434
rect 4318 17382 4328 17434
rect 4352 17382 4382 17434
rect 4382 17382 4394 17434
rect 4394 17382 4408 17434
rect 4432 17382 4446 17434
rect 4446 17382 4458 17434
rect 4458 17382 4488 17434
rect 4512 17382 4522 17434
rect 4522 17382 4568 17434
rect 4272 17380 4328 17382
rect 4352 17380 4408 17382
rect 4432 17380 4488 17382
rect 4512 17380 4568 17382
rect 4272 16346 4328 16348
rect 4352 16346 4408 16348
rect 4432 16346 4488 16348
rect 4512 16346 4568 16348
rect 4272 16294 4318 16346
rect 4318 16294 4328 16346
rect 4352 16294 4382 16346
rect 4382 16294 4394 16346
rect 4394 16294 4408 16346
rect 4432 16294 4446 16346
rect 4446 16294 4458 16346
rect 4458 16294 4488 16346
rect 4512 16294 4522 16346
rect 4522 16294 4568 16346
rect 4272 16292 4328 16294
rect 4352 16292 4408 16294
rect 4432 16292 4488 16294
rect 4512 16292 4568 16294
rect 3612 15802 3668 15804
rect 3692 15802 3748 15804
rect 3772 15802 3828 15804
rect 3852 15802 3908 15804
rect 3612 15750 3658 15802
rect 3658 15750 3668 15802
rect 3692 15750 3722 15802
rect 3722 15750 3734 15802
rect 3734 15750 3748 15802
rect 3772 15750 3786 15802
rect 3786 15750 3798 15802
rect 3798 15750 3828 15802
rect 3852 15750 3862 15802
rect 3862 15750 3908 15802
rect 3612 15748 3668 15750
rect 3692 15748 3748 15750
rect 3772 15748 3828 15750
rect 3852 15748 3908 15750
rect 4272 15258 4328 15260
rect 4352 15258 4408 15260
rect 4432 15258 4488 15260
rect 4512 15258 4568 15260
rect 4272 15206 4318 15258
rect 4318 15206 4328 15258
rect 4352 15206 4382 15258
rect 4382 15206 4394 15258
rect 4394 15206 4408 15258
rect 4432 15206 4446 15258
rect 4446 15206 4458 15258
rect 4458 15206 4488 15258
rect 4512 15206 4522 15258
rect 4522 15206 4568 15258
rect 4272 15204 4328 15206
rect 4352 15204 4408 15206
rect 4432 15204 4488 15206
rect 4512 15204 4568 15206
rect 3612 14714 3668 14716
rect 3692 14714 3748 14716
rect 3772 14714 3828 14716
rect 3852 14714 3908 14716
rect 3612 14662 3658 14714
rect 3658 14662 3668 14714
rect 3692 14662 3722 14714
rect 3722 14662 3734 14714
rect 3734 14662 3748 14714
rect 3772 14662 3786 14714
rect 3786 14662 3798 14714
rect 3798 14662 3828 14714
rect 3852 14662 3862 14714
rect 3862 14662 3908 14714
rect 3612 14660 3668 14662
rect 3692 14660 3748 14662
rect 3772 14660 3828 14662
rect 3852 14660 3908 14662
rect 4272 14170 4328 14172
rect 4352 14170 4408 14172
rect 4432 14170 4488 14172
rect 4512 14170 4568 14172
rect 4272 14118 4318 14170
rect 4318 14118 4328 14170
rect 4352 14118 4382 14170
rect 4382 14118 4394 14170
rect 4394 14118 4408 14170
rect 4432 14118 4446 14170
rect 4446 14118 4458 14170
rect 4458 14118 4488 14170
rect 4512 14118 4522 14170
rect 4522 14118 4568 14170
rect 4272 14116 4328 14118
rect 4352 14116 4408 14118
rect 4432 14116 4488 14118
rect 4512 14116 4568 14118
rect 3612 13626 3668 13628
rect 3692 13626 3748 13628
rect 3772 13626 3828 13628
rect 3852 13626 3908 13628
rect 3612 13574 3658 13626
rect 3658 13574 3668 13626
rect 3692 13574 3722 13626
rect 3722 13574 3734 13626
rect 3734 13574 3748 13626
rect 3772 13574 3786 13626
rect 3786 13574 3798 13626
rect 3798 13574 3828 13626
rect 3852 13574 3862 13626
rect 3862 13574 3908 13626
rect 3612 13572 3668 13574
rect 3692 13572 3748 13574
rect 3772 13572 3828 13574
rect 3852 13572 3908 13574
rect 4272 13082 4328 13084
rect 4352 13082 4408 13084
rect 4432 13082 4488 13084
rect 4512 13082 4568 13084
rect 4272 13030 4318 13082
rect 4318 13030 4328 13082
rect 4352 13030 4382 13082
rect 4382 13030 4394 13082
rect 4394 13030 4408 13082
rect 4432 13030 4446 13082
rect 4446 13030 4458 13082
rect 4458 13030 4488 13082
rect 4512 13030 4522 13082
rect 4522 13030 4568 13082
rect 4272 13028 4328 13030
rect 4352 13028 4408 13030
rect 4432 13028 4488 13030
rect 4512 13028 4568 13030
rect 3612 12538 3668 12540
rect 3692 12538 3748 12540
rect 3772 12538 3828 12540
rect 3852 12538 3908 12540
rect 3612 12486 3658 12538
rect 3658 12486 3668 12538
rect 3692 12486 3722 12538
rect 3722 12486 3734 12538
rect 3734 12486 3748 12538
rect 3772 12486 3786 12538
rect 3786 12486 3798 12538
rect 3798 12486 3828 12538
rect 3852 12486 3862 12538
rect 3862 12486 3908 12538
rect 3612 12484 3668 12486
rect 3692 12484 3748 12486
rect 3772 12484 3828 12486
rect 3852 12484 3908 12486
rect 4272 11994 4328 11996
rect 4352 11994 4408 11996
rect 4432 11994 4488 11996
rect 4512 11994 4568 11996
rect 4272 11942 4318 11994
rect 4318 11942 4328 11994
rect 4352 11942 4382 11994
rect 4382 11942 4394 11994
rect 4394 11942 4408 11994
rect 4432 11942 4446 11994
rect 4446 11942 4458 11994
rect 4458 11942 4488 11994
rect 4512 11942 4522 11994
rect 4522 11942 4568 11994
rect 4272 11940 4328 11942
rect 4352 11940 4408 11942
rect 4432 11940 4488 11942
rect 4512 11940 4568 11942
rect 3612 11450 3668 11452
rect 3692 11450 3748 11452
rect 3772 11450 3828 11452
rect 3852 11450 3908 11452
rect 3612 11398 3658 11450
rect 3658 11398 3668 11450
rect 3692 11398 3722 11450
rect 3722 11398 3734 11450
rect 3734 11398 3748 11450
rect 3772 11398 3786 11450
rect 3786 11398 3798 11450
rect 3798 11398 3828 11450
rect 3852 11398 3862 11450
rect 3862 11398 3908 11450
rect 3612 11396 3668 11398
rect 3692 11396 3748 11398
rect 3772 11396 3828 11398
rect 3852 11396 3908 11398
rect 3612 10362 3668 10364
rect 3692 10362 3748 10364
rect 3772 10362 3828 10364
rect 3852 10362 3908 10364
rect 3612 10310 3658 10362
rect 3658 10310 3668 10362
rect 3692 10310 3722 10362
rect 3722 10310 3734 10362
rect 3734 10310 3748 10362
rect 3772 10310 3786 10362
rect 3786 10310 3798 10362
rect 3798 10310 3828 10362
rect 3852 10310 3862 10362
rect 3862 10310 3908 10362
rect 3612 10308 3668 10310
rect 3692 10308 3748 10310
rect 3772 10308 3828 10310
rect 3852 10308 3908 10310
rect 4272 10906 4328 10908
rect 4352 10906 4408 10908
rect 4432 10906 4488 10908
rect 4512 10906 4568 10908
rect 4272 10854 4318 10906
rect 4318 10854 4328 10906
rect 4352 10854 4382 10906
rect 4382 10854 4394 10906
rect 4394 10854 4408 10906
rect 4432 10854 4446 10906
rect 4446 10854 4458 10906
rect 4458 10854 4488 10906
rect 4512 10854 4522 10906
rect 4522 10854 4568 10906
rect 4272 10852 4328 10854
rect 4352 10852 4408 10854
rect 4432 10852 4488 10854
rect 4512 10852 4568 10854
rect 846 7404 902 7440
rect 846 7384 848 7404
rect 848 7384 900 7404
rect 900 7384 902 7404
rect 4272 9818 4328 9820
rect 4352 9818 4408 9820
rect 4432 9818 4488 9820
rect 4512 9818 4568 9820
rect 4272 9766 4318 9818
rect 4318 9766 4328 9818
rect 4352 9766 4382 9818
rect 4382 9766 4394 9818
rect 4394 9766 4408 9818
rect 4432 9766 4446 9818
rect 4446 9766 4458 9818
rect 4458 9766 4488 9818
rect 4512 9766 4522 9818
rect 4522 9766 4568 9818
rect 4272 9764 4328 9766
rect 4352 9764 4408 9766
rect 4432 9764 4488 9766
rect 4512 9764 4568 9766
rect 3612 9274 3668 9276
rect 3692 9274 3748 9276
rect 3772 9274 3828 9276
rect 3852 9274 3908 9276
rect 3612 9222 3658 9274
rect 3658 9222 3668 9274
rect 3692 9222 3722 9274
rect 3722 9222 3734 9274
rect 3734 9222 3748 9274
rect 3772 9222 3786 9274
rect 3786 9222 3798 9274
rect 3798 9222 3828 9274
rect 3852 9222 3862 9274
rect 3862 9222 3908 9274
rect 3612 9220 3668 9222
rect 3692 9220 3748 9222
rect 3772 9220 3828 9222
rect 3852 9220 3908 9222
rect 4272 8730 4328 8732
rect 4352 8730 4408 8732
rect 4432 8730 4488 8732
rect 4512 8730 4568 8732
rect 4272 8678 4318 8730
rect 4318 8678 4328 8730
rect 4352 8678 4382 8730
rect 4382 8678 4394 8730
rect 4394 8678 4408 8730
rect 4432 8678 4446 8730
rect 4446 8678 4458 8730
rect 4458 8678 4488 8730
rect 4512 8678 4522 8730
rect 4522 8678 4568 8730
rect 4272 8676 4328 8678
rect 4352 8676 4408 8678
rect 4432 8676 4488 8678
rect 4512 8676 4568 8678
rect 1674 6840 1730 6896
rect 3612 8186 3668 8188
rect 3692 8186 3748 8188
rect 3772 8186 3828 8188
rect 3852 8186 3908 8188
rect 3612 8134 3658 8186
rect 3658 8134 3668 8186
rect 3692 8134 3722 8186
rect 3722 8134 3734 8186
rect 3734 8134 3748 8186
rect 3772 8134 3786 8186
rect 3786 8134 3798 8186
rect 3798 8134 3828 8186
rect 3852 8134 3862 8186
rect 3862 8134 3908 8186
rect 3612 8132 3668 8134
rect 3692 8132 3748 8134
rect 3772 8132 3828 8134
rect 3852 8132 3908 8134
rect 4272 7642 4328 7644
rect 4352 7642 4408 7644
rect 4432 7642 4488 7644
rect 4512 7642 4568 7644
rect 4272 7590 4318 7642
rect 4318 7590 4328 7642
rect 4352 7590 4382 7642
rect 4382 7590 4394 7642
rect 4394 7590 4408 7642
rect 4432 7590 4446 7642
rect 4446 7590 4458 7642
rect 4458 7590 4488 7642
rect 4512 7590 4522 7642
rect 4522 7590 4568 7642
rect 4272 7588 4328 7590
rect 4352 7588 4408 7590
rect 4432 7588 4488 7590
rect 4512 7588 4568 7590
rect 3612 7098 3668 7100
rect 3692 7098 3748 7100
rect 3772 7098 3828 7100
rect 3852 7098 3908 7100
rect 3612 7046 3658 7098
rect 3658 7046 3668 7098
rect 3692 7046 3722 7098
rect 3722 7046 3734 7098
rect 3734 7046 3748 7098
rect 3772 7046 3786 7098
rect 3786 7046 3798 7098
rect 3798 7046 3828 7098
rect 3852 7046 3862 7098
rect 3862 7046 3908 7098
rect 3612 7044 3668 7046
rect 3692 7044 3748 7046
rect 3772 7044 3828 7046
rect 3852 7044 3908 7046
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 4272 6554 4328 6556
rect 4352 6554 4408 6556
rect 4432 6554 4488 6556
rect 4512 6554 4568 6556
rect 4272 6502 4318 6554
rect 4318 6502 4328 6554
rect 4352 6502 4382 6554
rect 4382 6502 4394 6554
rect 4394 6502 4408 6554
rect 4432 6502 4446 6554
rect 4446 6502 4458 6554
rect 4458 6502 4488 6554
rect 4512 6502 4522 6554
rect 4522 6502 4568 6554
rect 4272 6500 4328 6502
rect 4352 6500 4408 6502
rect 4432 6500 4488 6502
rect 4512 6500 4568 6502
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 3612 6010 3668 6012
rect 3692 6010 3748 6012
rect 3772 6010 3828 6012
rect 3852 6010 3908 6012
rect 3612 5958 3658 6010
rect 3658 5958 3668 6010
rect 3692 5958 3722 6010
rect 3722 5958 3734 6010
rect 3734 5958 3748 6010
rect 3772 5958 3786 6010
rect 3786 5958 3798 6010
rect 3798 5958 3828 6010
rect 3852 5958 3862 6010
rect 3862 5958 3908 6010
rect 3612 5956 3668 5958
rect 3692 5956 3748 5958
rect 3772 5956 3828 5958
rect 3852 5956 3908 5958
rect 9585 22874 9641 22876
rect 9665 22874 9721 22876
rect 9745 22874 9801 22876
rect 9825 22874 9881 22876
rect 9585 22822 9631 22874
rect 9631 22822 9641 22874
rect 9665 22822 9695 22874
rect 9695 22822 9707 22874
rect 9707 22822 9721 22874
rect 9745 22822 9759 22874
rect 9759 22822 9771 22874
rect 9771 22822 9801 22874
rect 9825 22822 9835 22874
rect 9835 22822 9881 22874
rect 9585 22820 9641 22822
rect 9665 22820 9721 22822
rect 9745 22820 9801 22822
rect 9825 22820 9881 22822
rect 8925 22330 8981 22332
rect 9005 22330 9061 22332
rect 9085 22330 9141 22332
rect 9165 22330 9221 22332
rect 8925 22278 8971 22330
rect 8971 22278 8981 22330
rect 9005 22278 9035 22330
rect 9035 22278 9047 22330
rect 9047 22278 9061 22330
rect 9085 22278 9099 22330
rect 9099 22278 9111 22330
rect 9111 22278 9141 22330
rect 9165 22278 9175 22330
rect 9175 22278 9221 22330
rect 8925 22276 8981 22278
rect 9005 22276 9061 22278
rect 9085 22276 9141 22278
rect 9165 22276 9221 22278
rect 9585 21786 9641 21788
rect 9665 21786 9721 21788
rect 9745 21786 9801 21788
rect 9825 21786 9881 21788
rect 9585 21734 9631 21786
rect 9631 21734 9641 21786
rect 9665 21734 9695 21786
rect 9695 21734 9707 21786
rect 9707 21734 9721 21786
rect 9745 21734 9759 21786
rect 9759 21734 9771 21786
rect 9771 21734 9801 21786
rect 9825 21734 9835 21786
rect 9835 21734 9881 21786
rect 9585 21732 9641 21734
rect 9665 21732 9721 21734
rect 9745 21732 9801 21734
rect 9825 21732 9881 21734
rect 8925 21242 8981 21244
rect 9005 21242 9061 21244
rect 9085 21242 9141 21244
rect 9165 21242 9221 21244
rect 8925 21190 8971 21242
rect 8971 21190 8981 21242
rect 9005 21190 9035 21242
rect 9035 21190 9047 21242
rect 9047 21190 9061 21242
rect 9085 21190 9099 21242
rect 9099 21190 9111 21242
rect 9111 21190 9141 21242
rect 9165 21190 9175 21242
rect 9175 21190 9221 21242
rect 8925 21188 8981 21190
rect 9005 21188 9061 21190
rect 9085 21188 9141 21190
rect 9165 21188 9221 21190
rect 9585 20698 9641 20700
rect 9665 20698 9721 20700
rect 9745 20698 9801 20700
rect 9825 20698 9881 20700
rect 9585 20646 9631 20698
rect 9631 20646 9641 20698
rect 9665 20646 9695 20698
rect 9695 20646 9707 20698
rect 9707 20646 9721 20698
rect 9745 20646 9759 20698
rect 9759 20646 9771 20698
rect 9771 20646 9801 20698
rect 9825 20646 9835 20698
rect 9835 20646 9881 20698
rect 9585 20644 9641 20646
rect 9665 20644 9721 20646
rect 9745 20644 9801 20646
rect 9825 20644 9881 20646
rect 8925 20154 8981 20156
rect 9005 20154 9061 20156
rect 9085 20154 9141 20156
rect 9165 20154 9221 20156
rect 8925 20102 8971 20154
rect 8971 20102 8981 20154
rect 9005 20102 9035 20154
rect 9035 20102 9047 20154
rect 9047 20102 9061 20154
rect 9085 20102 9099 20154
rect 9099 20102 9111 20154
rect 9111 20102 9141 20154
rect 9165 20102 9175 20154
rect 9175 20102 9221 20154
rect 8925 20100 8981 20102
rect 9005 20100 9061 20102
rect 9085 20100 9141 20102
rect 9165 20100 9221 20102
rect 9585 19610 9641 19612
rect 9665 19610 9721 19612
rect 9745 19610 9801 19612
rect 9825 19610 9881 19612
rect 9585 19558 9631 19610
rect 9631 19558 9641 19610
rect 9665 19558 9695 19610
rect 9695 19558 9707 19610
rect 9707 19558 9721 19610
rect 9745 19558 9759 19610
rect 9759 19558 9771 19610
rect 9771 19558 9801 19610
rect 9825 19558 9835 19610
rect 9835 19558 9881 19610
rect 9585 19556 9641 19558
rect 9665 19556 9721 19558
rect 9745 19556 9801 19558
rect 9825 19556 9881 19558
rect 8925 19066 8981 19068
rect 9005 19066 9061 19068
rect 9085 19066 9141 19068
rect 9165 19066 9221 19068
rect 8925 19014 8971 19066
rect 8971 19014 8981 19066
rect 9005 19014 9035 19066
rect 9035 19014 9047 19066
rect 9047 19014 9061 19066
rect 9085 19014 9099 19066
rect 9099 19014 9111 19066
rect 9111 19014 9141 19066
rect 9165 19014 9175 19066
rect 9175 19014 9221 19066
rect 8925 19012 8981 19014
rect 9005 19012 9061 19014
rect 9085 19012 9141 19014
rect 9165 19012 9221 19014
rect 9585 18522 9641 18524
rect 9665 18522 9721 18524
rect 9745 18522 9801 18524
rect 9825 18522 9881 18524
rect 9585 18470 9631 18522
rect 9631 18470 9641 18522
rect 9665 18470 9695 18522
rect 9695 18470 9707 18522
rect 9707 18470 9721 18522
rect 9745 18470 9759 18522
rect 9759 18470 9771 18522
rect 9771 18470 9801 18522
rect 9825 18470 9835 18522
rect 9835 18470 9881 18522
rect 9585 18468 9641 18470
rect 9665 18468 9721 18470
rect 9745 18468 9801 18470
rect 9825 18468 9881 18470
rect 8925 17978 8981 17980
rect 9005 17978 9061 17980
rect 9085 17978 9141 17980
rect 9165 17978 9221 17980
rect 8925 17926 8971 17978
rect 8971 17926 8981 17978
rect 9005 17926 9035 17978
rect 9035 17926 9047 17978
rect 9047 17926 9061 17978
rect 9085 17926 9099 17978
rect 9099 17926 9111 17978
rect 9111 17926 9141 17978
rect 9165 17926 9175 17978
rect 9175 17926 9221 17978
rect 8925 17924 8981 17926
rect 9005 17924 9061 17926
rect 9085 17924 9141 17926
rect 9165 17924 9221 17926
rect 9585 17434 9641 17436
rect 9665 17434 9721 17436
rect 9745 17434 9801 17436
rect 9825 17434 9881 17436
rect 9585 17382 9631 17434
rect 9631 17382 9641 17434
rect 9665 17382 9695 17434
rect 9695 17382 9707 17434
rect 9707 17382 9721 17434
rect 9745 17382 9759 17434
rect 9759 17382 9771 17434
rect 9771 17382 9801 17434
rect 9825 17382 9835 17434
rect 9835 17382 9881 17434
rect 9585 17380 9641 17382
rect 9665 17380 9721 17382
rect 9745 17380 9801 17382
rect 9825 17380 9881 17382
rect 8925 16890 8981 16892
rect 9005 16890 9061 16892
rect 9085 16890 9141 16892
rect 9165 16890 9221 16892
rect 8925 16838 8971 16890
rect 8971 16838 8981 16890
rect 9005 16838 9035 16890
rect 9035 16838 9047 16890
rect 9047 16838 9061 16890
rect 9085 16838 9099 16890
rect 9099 16838 9111 16890
rect 9111 16838 9141 16890
rect 9165 16838 9175 16890
rect 9175 16838 9221 16890
rect 8925 16836 8981 16838
rect 9005 16836 9061 16838
rect 9085 16836 9141 16838
rect 9165 16836 9221 16838
rect 9585 16346 9641 16348
rect 9665 16346 9721 16348
rect 9745 16346 9801 16348
rect 9825 16346 9881 16348
rect 9585 16294 9631 16346
rect 9631 16294 9641 16346
rect 9665 16294 9695 16346
rect 9695 16294 9707 16346
rect 9707 16294 9721 16346
rect 9745 16294 9759 16346
rect 9759 16294 9771 16346
rect 9771 16294 9801 16346
rect 9825 16294 9835 16346
rect 9835 16294 9881 16346
rect 9585 16292 9641 16294
rect 9665 16292 9721 16294
rect 9745 16292 9801 16294
rect 9825 16292 9881 16294
rect 8925 15802 8981 15804
rect 9005 15802 9061 15804
rect 9085 15802 9141 15804
rect 9165 15802 9221 15804
rect 8925 15750 8971 15802
rect 8971 15750 8981 15802
rect 9005 15750 9035 15802
rect 9035 15750 9047 15802
rect 9047 15750 9061 15802
rect 9085 15750 9099 15802
rect 9099 15750 9111 15802
rect 9111 15750 9141 15802
rect 9165 15750 9175 15802
rect 9175 15750 9221 15802
rect 8925 15748 8981 15750
rect 9005 15748 9061 15750
rect 9085 15748 9141 15750
rect 9165 15748 9221 15750
rect 9585 15258 9641 15260
rect 9665 15258 9721 15260
rect 9745 15258 9801 15260
rect 9825 15258 9881 15260
rect 9585 15206 9631 15258
rect 9631 15206 9641 15258
rect 9665 15206 9695 15258
rect 9695 15206 9707 15258
rect 9707 15206 9721 15258
rect 9745 15206 9759 15258
rect 9759 15206 9771 15258
rect 9771 15206 9801 15258
rect 9825 15206 9835 15258
rect 9835 15206 9881 15258
rect 9585 15204 9641 15206
rect 9665 15204 9721 15206
rect 9745 15204 9801 15206
rect 9825 15204 9881 15206
rect 8925 14714 8981 14716
rect 9005 14714 9061 14716
rect 9085 14714 9141 14716
rect 9165 14714 9221 14716
rect 8925 14662 8971 14714
rect 8971 14662 8981 14714
rect 9005 14662 9035 14714
rect 9035 14662 9047 14714
rect 9047 14662 9061 14714
rect 9085 14662 9099 14714
rect 9099 14662 9111 14714
rect 9111 14662 9141 14714
rect 9165 14662 9175 14714
rect 9175 14662 9221 14714
rect 8925 14660 8981 14662
rect 9005 14660 9061 14662
rect 9085 14660 9141 14662
rect 9165 14660 9221 14662
rect 8925 13626 8981 13628
rect 9005 13626 9061 13628
rect 9085 13626 9141 13628
rect 9165 13626 9221 13628
rect 8925 13574 8971 13626
rect 8971 13574 8981 13626
rect 9005 13574 9035 13626
rect 9035 13574 9047 13626
rect 9047 13574 9061 13626
rect 9085 13574 9099 13626
rect 9099 13574 9111 13626
rect 9111 13574 9141 13626
rect 9165 13574 9175 13626
rect 9175 13574 9221 13626
rect 8925 13572 8981 13574
rect 9005 13572 9061 13574
rect 9085 13572 9141 13574
rect 9165 13572 9221 13574
rect 4272 5466 4328 5468
rect 4352 5466 4408 5468
rect 4432 5466 4488 5468
rect 4512 5466 4568 5468
rect 4272 5414 4318 5466
rect 4318 5414 4328 5466
rect 4352 5414 4382 5466
rect 4382 5414 4394 5466
rect 4394 5414 4408 5466
rect 4432 5414 4446 5466
rect 4446 5414 4458 5466
rect 4458 5414 4488 5466
rect 4512 5414 4522 5466
rect 4522 5414 4568 5466
rect 4272 5412 4328 5414
rect 4352 5412 4408 5414
rect 4432 5412 4488 5414
rect 4512 5412 4568 5414
rect 846 4936 902 4992
rect 3612 4922 3668 4924
rect 3692 4922 3748 4924
rect 3772 4922 3828 4924
rect 3852 4922 3908 4924
rect 3612 4870 3658 4922
rect 3658 4870 3668 4922
rect 3692 4870 3722 4922
rect 3722 4870 3734 4922
rect 3734 4870 3748 4922
rect 3772 4870 3786 4922
rect 3786 4870 3798 4922
rect 3798 4870 3828 4922
rect 3852 4870 3862 4922
rect 3862 4870 3908 4922
rect 3612 4868 3668 4870
rect 3692 4868 3748 4870
rect 3772 4868 3828 4870
rect 3852 4868 3908 4870
rect 846 4256 902 4312
rect 4272 4378 4328 4380
rect 4352 4378 4408 4380
rect 4432 4378 4488 4380
rect 4512 4378 4568 4380
rect 4272 4326 4318 4378
rect 4318 4326 4328 4378
rect 4352 4326 4382 4378
rect 4382 4326 4394 4378
rect 4394 4326 4408 4378
rect 4432 4326 4446 4378
rect 4446 4326 4458 4378
rect 4458 4326 4488 4378
rect 4512 4326 4522 4378
rect 4522 4326 4568 4378
rect 4272 4324 4328 4326
rect 4352 4324 4408 4326
rect 4432 4324 4488 4326
rect 4512 4324 4568 4326
rect 8925 12538 8981 12540
rect 9005 12538 9061 12540
rect 9085 12538 9141 12540
rect 9165 12538 9221 12540
rect 8925 12486 8971 12538
rect 8971 12486 8981 12538
rect 9005 12486 9035 12538
rect 9035 12486 9047 12538
rect 9047 12486 9061 12538
rect 9085 12486 9099 12538
rect 9099 12486 9111 12538
rect 9111 12486 9141 12538
rect 9165 12486 9175 12538
rect 9175 12486 9221 12538
rect 8925 12484 8981 12486
rect 9005 12484 9061 12486
rect 9085 12484 9141 12486
rect 9165 12484 9221 12486
rect 9585 14170 9641 14172
rect 9665 14170 9721 14172
rect 9745 14170 9801 14172
rect 9825 14170 9881 14172
rect 9585 14118 9631 14170
rect 9631 14118 9641 14170
rect 9665 14118 9695 14170
rect 9695 14118 9707 14170
rect 9707 14118 9721 14170
rect 9745 14118 9759 14170
rect 9759 14118 9771 14170
rect 9771 14118 9801 14170
rect 9825 14118 9835 14170
rect 9835 14118 9881 14170
rect 9585 14116 9641 14118
rect 9665 14116 9721 14118
rect 9745 14116 9801 14118
rect 9825 14116 9881 14118
rect 14238 23418 14294 23420
rect 14318 23418 14374 23420
rect 14398 23418 14454 23420
rect 14478 23418 14534 23420
rect 14238 23366 14284 23418
rect 14284 23366 14294 23418
rect 14318 23366 14348 23418
rect 14348 23366 14360 23418
rect 14360 23366 14374 23418
rect 14398 23366 14412 23418
rect 14412 23366 14424 23418
rect 14424 23366 14454 23418
rect 14478 23366 14488 23418
rect 14488 23366 14534 23418
rect 14238 23364 14294 23366
rect 14318 23364 14374 23366
rect 14398 23364 14454 23366
rect 14478 23364 14534 23366
rect 19551 23418 19607 23420
rect 19631 23418 19687 23420
rect 19711 23418 19767 23420
rect 19791 23418 19847 23420
rect 19551 23366 19597 23418
rect 19597 23366 19607 23418
rect 19631 23366 19661 23418
rect 19661 23366 19673 23418
rect 19673 23366 19687 23418
rect 19711 23366 19725 23418
rect 19725 23366 19737 23418
rect 19737 23366 19767 23418
rect 19791 23366 19801 23418
rect 19801 23366 19847 23418
rect 19551 23364 19607 23366
rect 19631 23364 19687 23366
rect 19711 23364 19767 23366
rect 19791 23364 19847 23366
rect 9585 13082 9641 13084
rect 9665 13082 9721 13084
rect 9745 13082 9801 13084
rect 9825 13082 9881 13084
rect 9585 13030 9631 13082
rect 9631 13030 9641 13082
rect 9665 13030 9695 13082
rect 9695 13030 9707 13082
rect 9707 13030 9721 13082
rect 9745 13030 9759 13082
rect 9759 13030 9771 13082
rect 9771 13030 9801 13082
rect 9825 13030 9835 13082
rect 9835 13030 9881 13082
rect 9585 13028 9641 13030
rect 9665 13028 9721 13030
rect 9745 13028 9801 13030
rect 9825 13028 9881 13030
rect 9585 11994 9641 11996
rect 9665 11994 9721 11996
rect 9745 11994 9801 11996
rect 9825 11994 9881 11996
rect 9585 11942 9631 11994
rect 9631 11942 9641 11994
rect 9665 11942 9695 11994
rect 9695 11942 9707 11994
rect 9707 11942 9721 11994
rect 9745 11942 9759 11994
rect 9759 11942 9771 11994
rect 9771 11942 9801 11994
rect 9825 11942 9835 11994
rect 9835 11942 9881 11994
rect 9585 11940 9641 11942
rect 9665 11940 9721 11942
rect 9745 11940 9801 11942
rect 9825 11940 9881 11942
rect 8925 11450 8981 11452
rect 9005 11450 9061 11452
rect 9085 11450 9141 11452
rect 9165 11450 9221 11452
rect 8925 11398 8971 11450
rect 8971 11398 8981 11450
rect 9005 11398 9035 11450
rect 9035 11398 9047 11450
rect 9047 11398 9061 11450
rect 9085 11398 9099 11450
rect 9099 11398 9111 11450
rect 9111 11398 9141 11450
rect 9165 11398 9175 11450
rect 9175 11398 9221 11450
rect 8925 11396 8981 11398
rect 9005 11396 9061 11398
rect 9085 11396 9141 11398
rect 9165 11396 9221 11398
rect 9585 10906 9641 10908
rect 9665 10906 9721 10908
rect 9745 10906 9801 10908
rect 9825 10906 9881 10908
rect 9585 10854 9631 10906
rect 9631 10854 9641 10906
rect 9665 10854 9695 10906
rect 9695 10854 9707 10906
rect 9707 10854 9721 10906
rect 9745 10854 9759 10906
rect 9759 10854 9771 10906
rect 9771 10854 9801 10906
rect 9825 10854 9835 10906
rect 9835 10854 9881 10906
rect 9585 10852 9641 10854
rect 9665 10852 9721 10854
rect 9745 10852 9801 10854
rect 9825 10852 9881 10854
rect 8925 10362 8981 10364
rect 9005 10362 9061 10364
rect 9085 10362 9141 10364
rect 9165 10362 9221 10364
rect 8925 10310 8971 10362
rect 8971 10310 8981 10362
rect 9005 10310 9035 10362
rect 9035 10310 9047 10362
rect 9047 10310 9061 10362
rect 9085 10310 9099 10362
rect 9099 10310 9111 10362
rect 9111 10310 9141 10362
rect 9165 10310 9175 10362
rect 9175 10310 9221 10362
rect 8925 10308 8981 10310
rect 9005 10308 9061 10310
rect 9085 10308 9141 10310
rect 9165 10308 9221 10310
rect 8925 9274 8981 9276
rect 9005 9274 9061 9276
rect 9085 9274 9141 9276
rect 9165 9274 9221 9276
rect 8925 9222 8971 9274
rect 8971 9222 8981 9274
rect 9005 9222 9035 9274
rect 9035 9222 9047 9274
rect 9047 9222 9061 9274
rect 9085 9222 9099 9274
rect 9099 9222 9111 9274
rect 9111 9222 9141 9274
rect 9165 9222 9175 9274
rect 9175 9222 9221 9274
rect 8925 9220 8981 9222
rect 9005 9220 9061 9222
rect 9085 9220 9141 9222
rect 9165 9220 9221 9222
rect 9585 9818 9641 9820
rect 9665 9818 9721 9820
rect 9745 9818 9801 9820
rect 9825 9818 9881 9820
rect 9585 9766 9631 9818
rect 9631 9766 9641 9818
rect 9665 9766 9695 9818
rect 9695 9766 9707 9818
rect 9707 9766 9721 9818
rect 9745 9766 9759 9818
rect 9759 9766 9771 9818
rect 9771 9766 9801 9818
rect 9825 9766 9835 9818
rect 9835 9766 9881 9818
rect 9585 9764 9641 9766
rect 9665 9764 9721 9766
rect 9745 9764 9801 9766
rect 9825 9764 9881 9766
rect 9585 8730 9641 8732
rect 9665 8730 9721 8732
rect 9745 8730 9801 8732
rect 9825 8730 9881 8732
rect 9585 8678 9631 8730
rect 9631 8678 9641 8730
rect 9665 8678 9695 8730
rect 9695 8678 9707 8730
rect 9707 8678 9721 8730
rect 9745 8678 9759 8730
rect 9759 8678 9771 8730
rect 9771 8678 9801 8730
rect 9825 8678 9835 8730
rect 9835 8678 9881 8730
rect 9585 8676 9641 8678
rect 9665 8676 9721 8678
rect 9745 8676 9801 8678
rect 9825 8676 9881 8678
rect 3612 3834 3668 3836
rect 3692 3834 3748 3836
rect 3772 3834 3828 3836
rect 3852 3834 3908 3836
rect 3612 3782 3658 3834
rect 3658 3782 3668 3834
rect 3692 3782 3722 3834
rect 3722 3782 3734 3834
rect 3734 3782 3748 3834
rect 3772 3782 3786 3834
rect 3786 3782 3798 3834
rect 3798 3782 3828 3834
rect 3852 3782 3862 3834
rect 3862 3782 3908 3834
rect 3612 3780 3668 3782
rect 3692 3780 3748 3782
rect 3772 3780 3828 3782
rect 3852 3780 3908 3782
rect 846 3304 902 3360
rect 4272 3290 4328 3292
rect 4352 3290 4408 3292
rect 4432 3290 4488 3292
rect 4512 3290 4568 3292
rect 4272 3238 4318 3290
rect 4318 3238 4328 3290
rect 4352 3238 4382 3290
rect 4382 3238 4394 3290
rect 4394 3238 4408 3290
rect 4432 3238 4446 3290
rect 4446 3238 4458 3290
rect 4458 3238 4488 3290
rect 4512 3238 4522 3290
rect 4522 3238 4568 3290
rect 4272 3236 4328 3238
rect 4352 3236 4408 3238
rect 4432 3236 4488 3238
rect 4512 3236 4568 3238
rect 3612 2746 3668 2748
rect 3692 2746 3748 2748
rect 3772 2746 3828 2748
rect 3852 2746 3908 2748
rect 3612 2694 3658 2746
rect 3658 2694 3668 2746
rect 3692 2694 3722 2746
rect 3722 2694 3734 2746
rect 3734 2694 3748 2746
rect 3772 2694 3786 2746
rect 3786 2694 3798 2746
rect 3798 2694 3828 2746
rect 3852 2694 3862 2746
rect 3862 2694 3908 2746
rect 3612 2692 3668 2694
rect 3692 2692 3748 2694
rect 3772 2692 3828 2694
rect 3852 2692 3908 2694
rect 4272 2202 4328 2204
rect 4352 2202 4408 2204
rect 4432 2202 4488 2204
rect 4512 2202 4568 2204
rect 4272 2150 4318 2202
rect 4318 2150 4328 2202
rect 4352 2150 4382 2202
rect 4382 2150 4394 2202
rect 4394 2150 4408 2202
rect 4432 2150 4446 2202
rect 4446 2150 4458 2202
rect 4458 2150 4488 2202
rect 4512 2150 4522 2202
rect 4522 2150 4568 2202
rect 4272 2148 4328 2150
rect 4352 2148 4408 2150
rect 4432 2148 4488 2150
rect 4512 2148 4568 2150
rect 8925 8186 8981 8188
rect 9005 8186 9061 8188
rect 9085 8186 9141 8188
rect 9165 8186 9221 8188
rect 8925 8134 8971 8186
rect 8971 8134 8981 8186
rect 9005 8134 9035 8186
rect 9035 8134 9047 8186
rect 9047 8134 9061 8186
rect 9085 8134 9099 8186
rect 9099 8134 9111 8186
rect 9111 8134 9141 8186
rect 9165 8134 9175 8186
rect 9175 8134 9221 8186
rect 8925 8132 8981 8134
rect 9005 8132 9061 8134
rect 9085 8132 9141 8134
rect 9165 8132 9221 8134
rect 8925 7098 8981 7100
rect 9005 7098 9061 7100
rect 9085 7098 9141 7100
rect 9165 7098 9221 7100
rect 8925 7046 8971 7098
rect 8971 7046 8981 7098
rect 9005 7046 9035 7098
rect 9035 7046 9047 7098
rect 9047 7046 9061 7098
rect 9085 7046 9099 7098
rect 9099 7046 9111 7098
rect 9111 7046 9141 7098
rect 9165 7046 9175 7098
rect 9175 7046 9221 7098
rect 8925 7044 8981 7046
rect 9005 7044 9061 7046
rect 9085 7044 9141 7046
rect 9165 7044 9221 7046
rect 9585 7642 9641 7644
rect 9665 7642 9721 7644
rect 9745 7642 9801 7644
rect 9825 7642 9881 7644
rect 9585 7590 9631 7642
rect 9631 7590 9641 7642
rect 9665 7590 9695 7642
rect 9695 7590 9707 7642
rect 9707 7590 9721 7642
rect 9745 7590 9759 7642
rect 9759 7590 9771 7642
rect 9771 7590 9801 7642
rect 9825 7590 9835 7642
rect 9835 7590 9881 7642
rect 9585 7588 9641 7590
rect 9665 7588 9721 7590
rect 9745 7588 9801 7590
rect 9825 7588 9881 7590
rect 9585 6554 9641 6556
rect 9665 6554 9721 6556
rect 9745 6554 9801 6556
rect 9825 6554 9881 6556
rect 9585 6502 9631 6554
rect 9631 6502 9641 6554
rect 9665 6502 9695 6554
rect 9695 6502 9707 6554
rect 9707 6502 9721 6554
rect 9745 6502 9759 6554
rect 9759 6502 9771 6554
rect 9771 6502 9801 6554
rect 9825 6502 9835 6554
rect 9835 6502 9881 6554
rect 9585 6500 9641 6502
rect 9665 6500 9721 6502
rect 9745 6500 9801 6502
rect 9825 6500 9881 6502
rect 8925 6010 8981 6012
rect 9005 6010 9061 6012
rect 9085 6010 9141 6012
rect 9165 6010 9221 6012
rect 8925 5958 8971 6010
rect 8971 5958 8981 6010
rect 9005 5958 9035 6010
rect 9035 5958 9047 6010
rect 9047 5958 9061 6010
rect 9085 5958 9099 6010
rect 9099 5958 9111 6010
rect 9111 5958 9141 6010
rect 9165 5958 9175 6010
rect 9175 5958 9221 6010
rect 8925 5956 8981 5958
rect 9005 5956 9061 5958
rect 9085 5956 9141 5958
rect 9165 5956 9221 5958
rect 8925 4922 8981 4924
rect 9005 4922 9061 4924
rect 9085 4922 9141 4924
rect 9165 4922 9221 4924
rect 8925 4870 8971 4922
rect 8971 4870 8981 4922
rect 9005 4870 9035 4922
rect 9035 4870 9047 4922
rect 9047 4870 9061 4922
rect 9085 4870 9099 4922
rect 9099 4870 9111 4922
rect 9111 4870 9141 4922
rect 9165 4870 9175 4922
rect 9175 4870 9221 4922
rect 8925 4868 8981 4870
rect 9005 4868 9061 4870
rect 9085 4868 9141 4870
rect 9165 4868 9221 4870
rect 9585 5466 9641 5468
rect 9665 5466 9721 5468
rect 9745 5466 9801 5468
rect 9825 5466 9881 5468
rect 9585 5414 9631 5466
rect 9631 5414 9641 5466
rect 9665 5414 9695 5466
rect 9695 5414 9707 5466
rect 9707 5414 9721 5466
rect 9745 5414 9759 5466
rect 9759 5414 9771 5466
rect 9771 5414 9801 5466
rect 9825 5414 9835 5466
rect 9835 5414 9881 5466
rect 9585 5412 9641 5414
rect 9665 5412 9721 5414
rect 9745 5412 9801 5414
rect 9825 5412 9881 5414
rect 9585 4378 9641 4380
rect 9665 4378 9721 4380
rect 9745 4378 9801 4380
rect 9825 4378 9881 4380
rect 9585 4326 9631 4378
rect 9631 4326 9641 4378
rect 9665 4326 9695 4378
rect 9695 4326 9707 4378
rect 9707 4326 9721 4378
rect 9745 4326 9759 4378
rect 9759 4326 9771 4378
rect 9771 4326 9801 4378
rect 9825 4326 9835 4378
rect 9835 4326 9881 4378
rect 9585 4324 9641 4326
rect 9665 4324 9721 4326
rect 9745 4324 9801 4326
rect 9825 4324 9881 4326
rect 8925 3834 8981 3836
rect 9005 3834 9061 3836
rect 9085 3834 9141 3836
rect 9165 3834 9221 3836
rect 8925 3782 8971 3834
rect 8971 3782 8981 3834
rect 9005 3782 9035 3834
rect 9035 3782 9047 3834
rect 9047 3782 9061 3834
rect 9085 3782 9099 3834
rect 9099 3782 9111 3834
rect 9111 3782 9141 3834
rect 9165 3782 9175 3834
rect 9175 3782 9221 3834
rect 8925 3780 8981 3782
rect 9005 3780 9061 3782
rect 9085 3780 9141 3782
rect 9165 3780 9221 3782
rect 9585 3290 9641 3292
rect 9665 3290 9721 3292
rect 9745 3290 9801 3292
rect 9825 3290 9881 3292
rect 9585 3238 9631 3290
rect 9631 3238 9641 3290
rect 9665 3238 9695 3290
rect 9695 3238 9707 3290
rect 9707 3238 9721 3290
rect 9745 3238 9759 3290
rect 9759 3238 9771 3290
rect 9771 3238 9801 3290
rect 9825 3238 9835 3290
rect 9835 3238 9881 3290
rect 9585 3236 9641 3238
rect 9665 3236 9721 3238
rect 9745 3236 9801 3238
rect 9825 3236 9881 3238
rect 8925 2746 8981 2748
rect 9005 2746 9061 2748
rect 9085 2746 9141 2748
rect 9165 2746 9221 2748
rect 8925 2694 8971 2746
rect 8971 2694 8981 2746
rect 9005 2694 9035 2746
rect 9035 2694 9047 2746
rect 9047 2694 9061 2746
rect 9085 2694 9099 2746
rect 9099 2694 9111 2746
rect 9111 2694 9141 2746
rect 9165 2694 9175 2746
rect 9175 2694 9221 2746
rect 8925 2692 8981 2694
rect 9005 2692 9061 2694
rect 9085 2692 9141 2694
rect 9165 2692 9221 2694
rect 9585 2202 9641 2204
rect 9665 2202 9721 2204
rect 9745 2202 9801 2204
rect 9825 2202 9881 2204
rect 9585 2150 9631 2202
rect 9631 2150 9641 2202
rect 9665 2150 9695 2202
rect 9695 2150 9707 2202
rect 9707 2150 9721 2202
rect 9745 2150 9759 2202
rect 9759 2150 9771 2202
rect 9771 2150 9801 2202
rect 9825 2150 9835 2202
rect 9835 2150 9881 2202
rect 9585 2148 9641 2150
rect 9665 2148 9721 2150
rect 9745 2148 9801 2150
rect 9825 2148 9881 2150
rect 14238 22330 14294 22332
rect 14318 22330 14374 22332
rect 14398 22330 14454 22332
rect 14478 22330 14534 22332
rect 14238 22278 14284 22330
rect 14284 22278 14294 22330
rect 14318 22278 14348 22330
rect 14348 22278 14360 22330
rect 14360 22278 14374 22330
rect 14398 22278 14412 22330
rect 14412 22278 14424 22330
rect 14424 22278 14454 22330
rect 14478 22278 14488 22330
rect 14488 22278 14534 22330
rect 14238 22276 14294 22278
rect 14318 22276 14374 22278
rect 14398 22276 14454 22278
rect 14478 22276 14534 22278
rect 14238 21242 14294 21244
rect 14318 21242 14374 21244
rect 14398 21242 14454 21244
rect 14478 21242 14534 21244
rect 14238 21190 14284 21242
rect 14284 21190 14294 21242
rect 14318 21190 14348 21242
rect 14348 21190 14360 21242
rect 14360 21190 14374 21242
rect 14398 21190 14412 21242
rect 14412 21190 14424 21242
rect 14424 21190 14454 21242
rect 14478 21190 14488 21242
rect 14488 21190 14534 21242
rect 14238 21188 14294 21190
rect 14318 21188 14374 21190
rect 14398 21188 14454 21190
rect 14478 21188 14534 21190
rect 14238 20154 14294 20156
rect 14318 20154 14374 20156
rect 14398 20154 14454 20156
rect 14478 20154 14534 20156
rect 14238 20102 14284 20154
rect 14284 20102 14294 20154
rect 14318 20102 14348 20154
rect 14348 20102 14360 20154
rect 14360 20102 14374 20154
rect 14398 20102 14412 20154
rect 14412 20102 14424 20154
rect 14424 20102 14454 20154
rect 14478 20102 14488 20154
rect 14488 20102 14534 20154
rect 14238 20100 14294 20102
rect 14318 20100 14374 20102
rect 14398 20100 14454 20102
rect 14478 20100 14534 20102
rect 14238 19066 14294 19068
rect 14318 19066 14374 19068
rect 14398 19066 14454 19068
rect 14478 19066 14534 19068
rect 14238 19014 14284 19066
rect 14284 19014 14294 19066
rect 14318 19014 14348 19066
rect 14348 19014 14360 19066
rect 14360 19014 14374 19066
rect 14398 19014 14412 19066
rect 14412 19014 14424 19066
rect 14424 19014 14454 19066
rect 14478 19014 14488 19066
rect 14488 19014 14534 19066
rect 14238 19012 14294 19014
rect 14318 19012 14374 19014
rect 14398 19012 14454 19014
rect 14478 19012 14534 19014
rect 14238 17978 14294 17980
rect 14318 17978 14374 17980
rect 14398 17978 14454 17980
rect 14478 17978 14534 17980
rect 14238 17926 14284 17978
rect 14284 17926 14294 17978
rect 14318 17926 14348 17978
rect 14348 17926 14360 17978
rect 14360 17926 14374 17978
rect 14398 17926 14412 17978
rect 14412 17926 14424 17978
rect 14424 17926 14454 17978
rect 14478 17926 14488 17978
rect 14488 17926 14534 17978
rect 14238 17924 14294 17926
rect 14318 17924 14374 17926
rect 14398 17924 14454 17926
rect 14478 17924 14534 17926
rect 14238 16890 14294 16892
rect 14318 16890 14374 16892
rect 14398 16890 14454 16892
rect 14478 16890 14534 16892
rect 14238 16838 14284 16890
rect 14284 16838 14294 16890
rect 14318 16838 14348 16890
rect 14348 16838 14360 16890
rect 14360 16838 14374 16890
rect 14398 16838 14412 16890
rect 14412 16838 14424 16890
rect 14424 16838 14454 16890
rect 14478 16838 14488 16890
rect 14488 16838 14534 16890
rect 14238 16836 14294 16838
rect 14318 16836 14374 16838
rect 14398 16836 14454 16838
rect 14478 16836 14534 16838
rect 14898 22874 14954 22876
rect 14978 22874 15034 22876
rect 15058 22874 15114 22876
rect 15138 22874 15194 22876
rect 14898 22822 14944 22874
rect 14944 22822 14954 22874
rect 14978 22822 15008 22874
rect 15008 22822 15020 22874
rect 15020 22822 15034 22874
rect 15058 22822 15072 22874
rect 15072 22822 15084 22874
rect 15084 22822 15114 22874
rect 15138 22822 15148 22874
rect 15148 22822 15194 22874
rect 14898 22820 14954 22822
rect 14978 22820 15034 22822
rect 15058 22820 15114 22822
rect 15138 22820 15194 22822
rect 14898 21786 14954 21788
rect 14978 21786 15034 21788
rect 15058 21786 15114 21788
rect 15138 21786 15194 21788
rect 14898 21734 14944 21786
rect 14944 21734 14954 21786
rect 14978 21734 15008 21786
rect 15008 21734 15020 21786
rect 15020 21734 15034 21786
rect 15058 21734 15072 21786
rect 15072 21734 15084 21786
rect 15084 21734 15114 21786
rect 15138 21734 15148 21786
rect 15148 21734 15194 21786
rect 14898 21732 14954 21734
rect 14978 21732 15034 21734
rect 15058 21732 15114 21734
rect 15138 21732 15194 21734
rect 14898 20698 14954 20700
rect 14978 20698 15034 20700
rect 15058 20698 15114 20700
rect 15138 20698 15194 20700
rect 14898 20646 14944 20698
rect 14944 20646 14954 20698
rect 14978 20646 15008 20698
rect 15008 20646 15020 20698
rect 15020 20646 15034 20698
rect 15058 20646 15072 20698
rect 15072 20646 15084 20698
rect 15084 20646 15114 20698
rect 15138 20646 15148 20698
rect 15148 20646 15194 20698
rect 14898 20644 14954 20646
rect 14978 20644 15034 20646
rect 15058 20644 15114 20646
rect 15138 20644 15194 20646
rect 14898 19610 14954 19612
rect 14978 19610 15034 19612
rect 15058 19610 15114 19612
rect 15138 19610 15194 19612
rect 14898 19558 14944 19610
rect 14944 19558 14954 19610
rect 14978 19558 15008 19610
rect 15008 19558 15020 19610
rect 15020 19558 15034 19610
rect 15058 19558 15072 19610
rect 15072 19558 15084 19610
rect 15084 19558 15114 19610
rect 15138 19558 15148 19610
rect 15148 19558 15194 19610
rect 14898 19556 14954 19558
rect 14978 19556 15034 19558
rect 15058 19556 15114 19558
rect 15138 19556 15194 19558
rect 14898 18522 14954 18524
rect 14978 18522 15034 18524
rect 15058 18522 15114 18524
rect 15138 18522 15194 18524
rect 14898 18470 14944 18522
rect 14944 18470 14954 18522
rect 14978 18470 15008 18522
rect 15008 18470 15020 18522
rect 15020 18470 15034 18522
rect 15058 18470 15072 18522
rect 15072 18470 15084 18522
rect 15084 18470 15114 18522
rect 15138 18470 15148 18522
rect 15148 18470 15194 18522
rect 14898 18468 14954 18470
rect 14978 18468 15034 18470
rect 15058 18468 15114 18470
rect 15138 18468 15194 18470
rect 14898 17434 14954 17436
rect 14978 17434 15034 17436
rect 15058 17434 15114 17436
rect 15138 17434 15194 17436
rect 14898 17382 14944 17434
rect 14944 17382 14954 17434
rect 14978 17382 15008 17434
rect 15008 17382 15020 17434
rect 15020 17382 15034 17434
rect 15058 17382 15072 17434
rect 15072 17382 15084 17434
rect 15084 17382 15114 17434
rect 15138 17382 15148 17434
rect 15148 17382 15194 17434
rect 14898 17380 14954 17382
rect 14978 17380 15034 17382
rect 15058 17380 15114 17382
rect 15138 17380 15194 17382
rect 14898 16346 14954 16348
rect 14978 16346 15034 16348
rect 15058 16346 15114 16348
rect 15138 16346 15194 16348
rect 14898 16294 14944 16346
rect 14944 16294 14954 16346
rect 14978 16294 15008 16346
rect 15008 16294 15020 16346
rect 15020 16294 15034 16346
rect 15058 16294 15072 16346
rect 15072 16294 15084 16346
rect 15084 16294 15114 16346
rect 15138 16294 15148 16346
rect 15148 16294 15194 16346
rect 14898 16292 14954 16294
rect 14978 16292 15034 16294
rect 15058 16292 15114 16294
rect 15138 16292 15194 16294
rect 14238 15802 14294 15804
rect 14318 15802 14374 15804
rect 14398 15802 14454 15804
rect 14478 15802 14534 15804
rect 14238 15750 14284 15802
rect 14284 15750 14294 15802
rect 14318 15750 14348 15802
rect 14348 15750 14360 15802
rect 14360 15750 14374 15802
rect 14398 15750 14412 15802
rect 14412 15750 14424 15802
rect 14424 15750 14454 15802
rect 14478 15750 14488 15802
rect 14488 15750 14534 15802
rect 14238 15748 14294 15750
rect 14318 15748 14374 15750
rect 14398 15748 14454 15750
rect 14478 15748 14534 15750
rect 14898 15258 14954 15260
rect 14978 15258 15034 15260
rect 15058 15258 15114 15260
rect 15138 15258 15194 15260
rect 14898 15206 14944 15258
rect 14944 15206 14954 15258
rect 14978 15206 15008 15258
rect 15008 15206 15020 15258
rect 15020 15206 15034 15258
rect 15058 15206 15072 15258
rect 15072 15206 15084 15258
rect 15084 15206 15114 15258
rect 15138 15206 15148 15258
rect 15148 15206 15194 15258
rect 14898 15204 14954 15206
rect 14978 15204 15034 15206
rect 15058 15204 15114 15206
rect 15138 15204 15194 15206
rect 14238 14714 14294 14716
rect 14318 14714 14374 14716
rect 14398 14714 14454 14716
rect 14478 14714 14534 14716
rect 14238 14662 14284 14714
rect 14284 14662 14294 14714
rect 14318 14662 14348 14714
rect 14348 14662 14360 14714
rect 14360 14662 14374 14714
rect 14398 14662 14412 14714
rect 14412 14662 14424 14714
rect 14424 14662 14454 14714
rect 14478 14662 14488 14714
rect 14488 14662 14534 14714
rect 14238 14660 14294 14662
rect 14318 14660 14374 14662
rect 14398 14660 14454 14662
rect 14478 14660 14534 14662
rect 14898 14170 14954 14172
rect 14978 14170 15034 14172
rect 15058 14170 15114 14172
rect 15138 14170 15194 14172
rect 14898 14118 14944 14170
rect 14944 14118 14954 14170
rect 14978 14118 15008 14170
rect 15008 14118 15020 14170
rect 15020 14118 15034 14170
rect 15058 14118 15072 14170
rect 15072 14118 15084 14170
rect 15084 14118 15114 14170
rect 15138 14118 15148 14170
rect 15148 14118 15194 14170
rect 14898 14116 14954 14118
rect 14978 14116 15034 14118
rect 15058 14116 15114 14118
rect 15138 14116 15194 14118
rect 14238 13626 14294 13628
rect 14318 13626 14374 13628
rect 14398 13626 14454 13628
rect 14478 13626 14534 13628
rect 14238 13574 14284 13626
rect 14284 13574 14294 13626
rect 14318 13574 14348 13626
rect 14348 13574 14360 13626
rect 14360 13574 14374 13626
rect 14398 13574 14412 13626
rect 14412 13574 14424 13626
rect 14424 13574 14454 13626
rect 14478 13574 14488 13626
rect 14488 13574 14534 13626
rect 14238 13572 14294 13574
rect 14318 13572 14374 13574
rect 14398 13572 14454 13574
rect 14478 13572 14534 13574
rect 14898 13082 14954 13084
rect 14978 13082 15034 13084
rect 15058 13082 15114 13084
rect 15138 13082 15194 13084
rect 14898 13030 14944 13082
rect 14944 13030 14954 13082
rect 14978 13030 15008 13082
rect 15008 13030 15020 13082
rect 15020 13030 15034 13082
rect 15058 13030 15072 13082
rect 15072 13030 15084 13082
rect 15084 13030 15114 13082
rect 15138 13030 15148 13082
rect 15148 13030 15194 13082
rect 14898 13028 14954 13030
rect 14978 13028 15034 13030
rect 15058 13028 15114 13030
rect 15138 13028 15194 13030
rect 14238 12538 14294 12540
rect 14318 12538 14374 12540
rect 14398 12538 14454 12540
rect 14478 12538 14534 12540
rect 14238 12486 14284 12538
rect 14284 12486 14294 12538
rect 14318 12486 14348 12538
rect 14348 12486 14360 12538
rect 14360 12486 14374 12538
rect 14398 12486 14412 12538
rect 14412 12486 14424 12538
rect 14424 12486 14454 12538
rect 14478 12486 14488 12538
rect 14488 12486 14534 12538
rect 14238 12484 14294 12486
rect 14318 12484 14374 12486
rect 14398 12484 14454 12486
rect 14478 12484 14534 12486
rect 14898 11994 14954 11996
rect 14978 11994 15034 11996
rect 15058 11994 15114 11996
rect 15138 11994 15194 11996
rect 14898 11942 14944 11994
rect 14944 11942 14954 11994
rect 14978 11942 15008 11994
rect 15008 11942 15020 11994
rect 15020 11942 15034 11994
rect 15058 11942 15072 11994
rect 15072 11942 15084 11994
rect 15084 11942 15114 11994
rect 15138 11942 15148 11994
rect 15148 11942 15194 11994
rect 14898 11940 14954 11942
rect 14978 11940 15034 11942
rect 15058 11940 15114 11942
rect 15138 11940 15194 11942
rect 14238 11450 14294 11452
rect 14318 11450 14374 11452
rect 14398 11450 14454 11452
rect 14478 11450 14534 11452
rect 14238 11398 14284 11450
rect 14284 11398 14294 11450
rect 14318 11398 14348 11450
rect 14348 11398 14360 11450
rect 14360 11398 14374 11450
rect 14398 11398 14412 11450
rect 14412 11398 14424 11450
rect 14424 11398 14454 11450
rect 14478 11398 14488 11450
rect 14488 11398 14534 11450
rect 14238 11396 14294 11398
rect 14318 11396 14374 11398
rect 14398 11396 14454 11398
rect 14478 11396 14534 11398
rect 14898 10906 14954 10908
rect 14978 10906 15034 10908
rect 15058 10906 15114 10908
rect 15138 10906 15194 10908
rect 14898 10854 14944 10906
rect 14944 10854 14954 10906
rect 14978 10854 15008 10906
rect 15008 10854 15020 10906
rect 15020 10854 15034 10906
rect 15058 10854 15072 10906
rect 15072 10854 15084 10906
rect 15084 10854 15114 10906
rect 15138 10854 15148 10906
rect 15148 10854 15194 10906
rect 14898 10852 14954 10854
rect 14978 10852 15034 10854
rect 15058 10852 15114 10854
rect 15138 10852 15194 10854
rect 14238 10362 14294 10364
rect 14318 10362 14374 10364
rect 14398 10362 14454 10364
rect 14478 10362 14534 10364
rect 14238 10310 14284 10362
rect 14284 10310 14294 10362
rect 14318 10310 14348 10362
rect 14348 10310 14360 10362
rect 14360 10310 14374 10362
rect 14398 10310 14412 10362
rect 14412 10310 14424 10362
rect 14424 10310 14454 10362
rect 14478 10310 14488 10362
rect 14488 10310 14534 10362
rect 14238 10308 14294 10310
rect 14318 10308 14374 10310
rect 14398 10308 14454 10310
rect 14478 10308 14534 10310
rect 14238 9274 14294 9276
rect 14318 9274 14374 9276
rect 14398 9274 14454 9276
rect 14478 9274 14534 9276
rect 14238 9222 14284 9274
rect 14284 9222 14294 9274
rect 14318 9222 14348 9274
rect 14348 9222 14360 9274
rect 14360 9222 14374 9274
rect 14398 9222 14412 9274
rect 14412 9222 14424 9274
rect 14424 9222 14454 9274
rect 14478 9222 14488 9274
rect 14488 9222 14534 9274
rect 14238 9220 14294 9222
rect 14318 9220 14374 9222
rect 14398 9220 14454 9222
rect 14478 9220 14534 9222
rect 14238 8186 14294 8188
rect 14318 8186 14374 8188
rect 14398 8186 14454 8188
rect 14478 8186 14534 8188
rect 14238 8134 14284 8186
rect 14284 8134 14294 8186
rect 14318 8134 14348 8186
rect 14348 8134 14360 8186
rect 14360 8134 14374 8186
rect 14398 8134 14412 8186
rect 14412 8134 14424 8186
rect 14424 8134 14454 8186
rect 14478 8134 14488 8186
rect 14488 8134 14534 8186
rect 14238 8132 14294 8134
rect 14318 8132 14374 8134
rect 14398 8132 14454 8134
rect 14478 8132 14534 8134
rect 14898 9818 14954 9820
rect 14978 9818 15034 9820
rect 15058 9818 15114 9820
rect 15138 9818 15194 9820
rect 14898 9766 14944 9818
rect 14944 9766 14954 9818
rect 14978 9766 15008 9818
rect 15008 9766 15020 9818
rect 15020 9766 15034 9818
rect 15058 9766 15072 9818
rect 15072 9766 15084 9818
rect 15084 9766 15114 9818
rect 15138 9766 15148 9818
rect 15148 9766 15194 9818
rect 14898 9764 14954 9766
rect 14978 9764 15034 9766
rect 15058 9764 15114 9766
rect 15138 9764 15194 9766
rect 14238 7098 14294 7100
rect 14318 7098 14374 7100
rect 14398 7098 14454 7100
rect 14478 7098 14534 7100
rect 14238 7046 14284 7098
rect 14284 7046 14294 7098
rect 14318 7046 14348 7098
rect 14348 7046 14360 7098
rect 14360 7046 14374 7098
rect 14398 7046 14412 7098
rect 14412 7046 14424 7098
rect 14424 7046 14454 7098
rect 14478 7046 14488 7098
rect 14488 7046 14534 7098
rect 14238 7044 14294 7046
rect 14318 7044 14374 7046
rect 14398 7044 14454 7046
rect 14478 7044 14534 7046
rect 14898 8730 14954 8732
rect 14978 8730 15034 8732
rect 15058 8730 15114 8732
rect 15138 8730 15194 8732
rect 14898 8678 14944 8730
rect 14944 8678 14954 8730
rect 14978 8678 15008 8730
rect 15008 8678 15020 8730
rect 15020 8678 15034 8730
rect 15058 8678 15072 8730
rect 15072 8678 15084 8730
rect 15084 8678 15114 8730
rect 15138 8678 15148 8730
rect 15148 8678 15194 8730
rect 14898 8676 14954 8678
rect 14978 8676 15034 8678
rect 15058 8676 15114 8678
rect 15138 8676 15194 8678
rect 20211 22874 20267 22876
rect 20291 22874 20347 22876
rect 20371 22874 20427 22876
rect 20451 22874 20507 22876
rect 20211 22822 20257 22874
rect 20257 22822 20267 22874
rect 20291 22822 20321 22874
rect 20321 22822 20333 22874
rect 20333 22822 20347 22874
rect 20371 22822 20385 22874
rect 20385 22822 20397 22874
rect 20397 22822 20427 22874
rect 20451 22822 20461 22874
rect 20461 22822 20507 22874
rect 20211 22820 20267 22822
rect 20291 22820 20347 22822
rect 20371 22820 20427 22822
rect 20451 22820 20507 22822
rect 19551 22330 19607 22332
rect 19631 22330 19687 22332
rect 19711 22330 19767 22332
rect 19791 22330 19847 22332
rect 19551 22278 19597 22330
rect 19597 22278 19607 22330
rect 19631 22278 19661 22330
rect 19661 22278 19673 22330
rect 19673 22278 19687 22330
rect 19711 22278 19725 22330
rect 19725 22278 19737 22330
rect 19737 22278 19767 22330
rect 19791 22278 19801 22330
rect 19801 22278 19847 22330
rect 19551 22276 19607 22278
rect 19631 22276 19687 22278
rect 19711 22276 19767 22278
rect 19791 22276 19847 22278
rect 19551 21242 19607 21244
rect 19631 21242 19687 21244
rect 19711 21242 19767 21244
rect 19791 21242 19847 21244
rect 19551 21190 19597 21242
rect 19597 21190 19607 21242
rect 19631 21190 19661 21242
rect 19661 21190 19673 21242
rect 19673 21190 19687 21242
rect 19711 21190 19725 21242
rect 19725 21190 19737 21242
rect 19737 21190 19767 21242
rect 19791 21190 19801 21242
rect 19801 21190 19847 21242
rect 19551 21188 19607 21190
rect 19631 21188 19687 21190
rect 19711 21188 19767 21190
rect 19791 21188 19847 21190
rect 20211 21786 20267 21788
rect 20291 21786 20347 21788
rect 20371 21786 20427 21788
rect 20451 21786 20507 21788
rect 20211 21734 20257 21786
rect 20257 21734 20267 21786
rect 20291 21734 20321 21786
rect 20321 21734 20333 21786
rect 20333 21734 20347 21786
rect 20371 21734 20385 21786
rect 20385 21734 20397 21786
rect 20397 21734 20427 21786
rect 20451 21734 20461 21786
rect 20461 21734 20507 21786
rect 20211 21732 20267 21734
rect 20291 21732 20347 21734
rect 20371 21732 20427 21734
rect 20451 21732 20507 21734
rect 20211 20698 20267 20700
rect 20291 20698 20347 20700
rect 20371 20698 20427 20700
rect 20451 20698 20507 20700
rect 20211 20646 20257 20698
rect 20257 20646 20267 20698
rect 20291 20646 20321 20698
rect 20321 20646 20333 20698
rect 20333 20646 20347 20698
rect 20371 20646 20385 20698
rect 20385 20646 20397 20698
rect 20397 20646 20427 20698
rect 20451 20646 20461 20698
rect 20461 20646 20507 20698
rect 20211 20644 20267 20646
rect 20291 20644 20347 20646
rect 20371 20644 20427 20646
rect 20451 20644 20507 20646
rect 19551 20154 19607 20156
rect 19631 20154 19687 20156
rect 19711 20154 19767 20156
rect 19791 20154 19847 20156
rect 19551 20102 19597 20154
rect 19597 20102 19607 20154
rect 19631 20102 19661 20154
rect 19661 20102 19673 20154
rect 19673 20102 19687 20154
rect 19711 20102 19725 20154
rect 19725 20102 19737 20154
rect 19737 20102 19767 20154
rect 19791 20102 19801 20154
rect 19801 20102 19847 20154
rect 19551 20100 19607 20102
rect 19631 20100 19687 20102
rect 19711 20100 19767 20102
rect 19791 20100 19847 20102
rect 20211 19610 20267 19612
rect 20291 19610 20347 19612
rect 20371 19610 20427 19612
rect 20451 19610 20507 19612
rect 20211 19558 20257 19610
rect 20257 19558 20267 19610
rect 20291 19558 20321 19610
rect 20321 19558 20333 19610
rect 20333 19558 20347 19610
rect 20371 19558 20385 19610
rect 20385 19558 20397 19610
rect 20397 19558 20427 19610
rect 20451 19558 20461 19610
rect 20461 19558 20507 19610
rect 20211 19556 20267 19558
rect 20291 19556 20347 19558
rect 20371 19556 20427 19558
rect 20451 19556 20507 19558
rect 19551 19066 19607 19068
rect 19631 19066 19687 19068
rect 19711 19066 19767 19068
rect 19791 19066 19847 19068
rect 19551 19014 19597 19066
rect 19597 19014 19607 19066
rect 19631 19014 19661 19066
rect 19661 19014 19673 19066
rect 19673 19014 19687 19066
rect 19711 19014 19725 19066
rect 19725 19014 19737 19066
rect 19737 19014 19767 19066
rect 19791 19014 19801 19066
rect 19801 19014 19847 19066
rect 19551 19012 19607 19014
rect 19631 19012 19687 19014
rect 19711 19012 19767 19014
rect 19791 19012 19847 19014
rect 20211 18522 20267 18524
rect 20291 18522 20347 18524
rect 20371 18522 20427 18524
rect 20451 18522 20507 18524
rect 20211 18470 20257 18522
rect 20257 18470 20267 18522
rect 20291 18470 20321 18522
rect 20321 18470 20333 18522
rect 20333 18470 20347 18522
rect 20371 18470 20385 18522
rect 20385 18470 20397 18522
rect 20397 18470 20427 18522
rect 20451 18470 20461 18522
rect 20461 18470 20507 18522
rect 20211 18468 20267 18470
rect 20291 18468 20347 18470
rect 20371 18468 20427 18470
rect 20451 18468 20507 18470
rect 19551 17978 19607 17980
rect 19631 17978 19687 17980
rect 19711 17978 19767 17980
rect 19791 17978 19847 17980
rect 19551 17926 19597 17978
rect 19597 17926 19607 17978
rect 19631 17926 19661 17978
rect 19661 17926 19673 17978
rect 19673 17926 19687 17978
rect 19711 17926 19725 17978
rect 19725 17926 19737 17978
rect 19737 17926 19767 17978
rect 19791 17926 19801 17978
rect 19801 17926 19847 17978
rect 19551 17924 19607 17926
rect 19631 17924 19687 17926
rect 19711 17924 19767 17926
rect 19791 17924 19847 17926
rect 22006 20440 22062 20496
rect 20211 17434 20267 17436
rect 20291 17434 20347 17436
rect 20371 17434 20427 17436
rect 20451 17434 20507 17436
rect 20211 17382 20257 17434
rect 20257 17382 20267 17434
rect 20291 17382 20321 17434
rect 20321 17382 20333 17434
rect 20333 17382 20347 17434
rect 20371 17382 20385 17434
rect 20385 17382 20397 17434
rect 20397 17382 20427 17434
rect 20451 17382 20461 17434
rect 20461 17382 20507 17434
rect 20211 17380 20267 17382
rect 20291 17380 20347 17382
rect 20371 17380 20427 17382
rect 20451 17380 20507 17382
rect 19551 16890 19607 16892
rect 19631 16890 19687 16892
rect 19711 16890 19767 16892
rect 19791 16890 19847 16892
rect 19551 16838 19597 16890
rect 19597 16838 19607 16890
rect 19631 16838 19661 16890
rect 19661 16838 19673 16890
rect 19673 16838 19687 16890
rect 19711 16838 19725 16890
rect 19725 16838 19737 16890
rect 19737 16838 19767 16890
rect 19791 16838 19801 16890
rect 19801 16838 19847 16890
rect 19551 16836 19607 16838
rect 19631 16836 19687 16838
rect 19711 16836 19767 16838
rect 19791 16836 19847 16838
rect 20211 16346 20267 16348
rect 20291 16346 20347 16348
rect 20371 16346 20427 16348
rect 20451 16346 20507 16348
rect 20211 16294 20257 16346
rect 20257 16294 20267 16346
rect 20291 16294 20321 16346
rect 20321 16294 20333 16346
rect 20333 16294 20347 16346
rect 20371 16294 20385 16346
rect 20385 16294 20397 16346
rect 20397 16294 20427 16346
rect 20451 16294 20461 16346
rect 20461 16294 20507 16346
rect 20211 16292 20267 16294
rect 20291 16292 20347 16294
rect 20371 16292 20427 16294
rect 20451 16292 20507 16294
rect 19551 15802 19607 15804
rect 19631 15802 19687 15804
rect 19711 15802 19767 15804
rect 19791 15802 19847 15804
rect 19551 15750 19597 15802
rect 19597 15750 19607 15802
rect 19631 15750 19661 15802
rect 19661 15750 19673 15802
rect 19673 15750 19687 15802
rect 19711 15750 19725 15802
rect 19725 15750 19737 15802
rect 19737 15750 19767 15802
rect 19791 15750 19801 15802
rect 19801 15750 19847 15802
rect 19551 15748 19607 15750
rect 19631 15748 19687 15750
rect 19711 15748 19767 15750
rect 19791 15748 19847 15750
rect 20211 15258 20267 15260
rect 20291 15258 20347 15260
rect 20371 15258 20427 15260
rect 20451 15258 20507 15260
rect 20211 15206 20257 15258
rect 20257 15206 20267 15258
rect 20291 15206 20321 15258
rect 20321 15206 20333 15258
rect 20333 15206 20347 15258
rect 20371 15206 20385 15258
rect 20385 15206 20397 15258
rect 20397 15206 20427 15258
rect 20451 15206 20461 15258
rect 20461 15206 20507 15258
rect 20211 15204 20267 15206
rect 20291 15204 20347 15206
rect 20371 15204 20427 15206
rect 20451 15204 20507 15206
rect 22006 19796 22008 19816
rect 22008 19796 22060 19816
rect 22060 19796 22062 19816
rect 22006 19760 22062 19796
rect 19551 14714 19607 14716
rect 19631 14714 19687 14716
rect 19711 14714 19767 14716
rect 19791 14714 19847 14716
rect 19551 14662 19597 14714
rect 19597 14662 19607 14714
rect 19631 14662 19661 14714
rect 19661 14662 19673 14714
rect 19673 14662 19687 14714
rect 19711 14662 19725 14714
rect 19725 14662 19737 14714
rect 19737 14662 19767 14714
rect 19791 14662 19801 14714
rect 19801 14662 19847 14714
rect 19551 14660 19607 14662
rect 19631 14660 19687 14662
rect 19711 14660 19767 14662
rect 19791 14660 19847 14662
rect 14898 7642 14954 7644
rect 14978 7642 15034 7644
rect 15058 7642 15114 7644
rect 15138 7642 15194 7644
rect 14898 7590 14944 7642
rect 14944 7590 14954 7642
rect 14978 7590 15008 7642
rect 15008 7590 15020 7642
rect 15020 7590 15034 7642
rect 15058 7590 15072 7642
rect 15072 7590 15084 7642
rect 15084 7590 15114 7642
rect 15138 7590 15148 7642
rect 15148 7590 15194 7642
rect 14898 7588 14954 7590
rect 14978 7588 15034 7590
rect 15058 7588 15114 7590
rect 15138 7588 15194 7590
rect 14898 6554 14954 6556
rect 14978 6554 15034 6556
rect 15058 6554 15114 6556
rect 15138 6554 15194 6556
rect 14898 6502 14944 6554
rect 14944 6502 14954 6554
rect 14978 6502 15008 6554
rect 15008 6502 15020 6554
rect 15020 6502 15034 6554
rect 15058 6502 15072 6554
rect 15072 6502 15084 6554
rect 15084 6502 15114 6554
rect 15138 6502 15148 6554
rect 15148 6502 15194 6554
rect 14898 6500 14954 6502
rect 14978 6500 15034 6502
rect 15058 6500 15114 6502
rect 15138 6500 15194 6502
rect 14238 6010 14294 6012
rect 14318 6010 14374 6012
rect 14398 6010 14454 6012
rect 14478 6010 14534 6012
rect 14238 5958 14284 6010
rect 14284 5958 14294 6010
rect 14318 5958 14348 6010
rect 14348 5958 14360 6010
rect 14360 5958 14374 6010
rect 14398 5958 14412 6010
rect 14412 5958 14424 6010
rect 14424 5958 14454 6010
rect 14478 5958 14488 6010
rect 14488 5958 14534 6010
rect 14238 5956 14294 5958
rect 14318 5956 14374 5958
rect 14398 5956 14454 5958
rect 14478 5956 14534 5958
rect 14238 4922 14294 4924
rect 14318 4922 14374 4924
rect 14398 4922 14454 4924
rect 14478 4922 14534 4924
rect 14238 4870 14284 4922
rect 14284 4870 14294 4922
rect 14318 4870 14348 4922
rect 14348 4870 14360 4922
rect 14360 4870 14374 4922
rect 14398 4870 14412 4922
rect 14412 4870 14424 4922
rect 14424 4870 14454 4922
rect 14478 4870 14488 4922
rect 14488 4870 14534 4922
rect 14238 4868 14294 4870
rect 14318 4868 14374 4870
rect 14398 4868 14454 4870
rect 14478 4868 14534 4870
rect 14898 5466 14954 5468
rect 14978 5466 15034 5468
rect 15058 5466 15114 5468
rect 15138 5466 15194 5468
rect 14898 5414 14944 5466
rect 14944 5414 14954 5466
rect 14978 5414 15008 5466
rect 15008 5414 15020 5466
rect 15020 5414 15034 5466
rect 15058 5414 15072 5466
rect 15072 5414 15084 5466
rect 15084 5414 15114 5466
rect 15138 5414 15148 5466
rect 15148 5414 15194 5466
rect 14898 5412 14954 5414
rect 14978 5412 15034 5414
rect 15058 5412 15114 5414
rect 15138 5412 15194 5414
rect 14898 4378 14954 4380
rect 14978 4378 15034 4380
rect 15058 4378 15114 4380
rect 15138 4378 15194 4380
rect 14898 4326 14944 4378
rect 14944 4326 14954 4378
rect 14978 4326 15008 4378
rect 15008 4326 15020 4378
rect 15020 4326 15034 4378
rect 15058 4326 15072 4378
rect 15072 4326 15084 4378
rect 15084 4326 15114 4378
rect 15138 4326 15148 4378
rect 15148 4326 15194 4378
rect 14898 4324 14954 4326
rect 14978 4324 15034 4326
rect 15058 4324 15114 4326
rect 15138 4324 15194 4326
rect 14238 3834 14294 3836
rect 14318 3834 14374 3836
rect 14398 3834 14454 3836
rect 14478 3834 14534 3836
rect 14238 3782 14284 3834
rect 14284 3782 14294 3834
rect 14318 3782 14348 3834
rect 14348 3782 14360 3834
rect 14360 3782 14374 3834
rect 14398 3782 14412 3834
rect 14412 3782 14424 3834
rect 14424 3782 14454 3834
rect 14478 3782 14488 3834
rect 14488 3782 14534 3834
rect 14238 3780 14294 3782
rect 14318 3780 14374 3782
rect 14398 3780 14454 3782
rect 14478 3780 14534 3782
rect 14898 3290 14954 3292
rect 14978 3290 15034 3292
rect 15058 3290 15114 3292
rect 15138 3290 15194 3292
rect 14898 3238 14944 3290
rect 14944 3238 14954 3290
rect 14978 3238 15008 3290
rect 15008 3238 15020 3290
rect 15020 3238 15034 3290
rect 15058 3238 15072 3290
rect 15072 3238 15084 3290
rect 15084 3238 15114 3290
rect 15138 3238 15148 3290
rect 15148 3238 15194 3290
rect 14898 3236 14954 3238
rect 14978 3236 15034 3238
rect 15058 3236 15114 3238
rect 15138 3236 15194 3238
rect 14238 2746 14294 2748
rect 14318 2746 14374 2748
rect 14398 2746 14454 2748
rect 14478 2746 14534 2748
rect 14238 2694 14284 2746
rect 14284 2694 14294 2746
rect 14318 2694 14348 2746
rect 14348 2694 14360 2746
rect 14360 2694 14374 2746
rect 14398 2694 14412 2746
rect 14412 2694 14424 2746
rect 14424 2694 14454 2746
rect 14478 2694 14488 2746
rect 14488 2694 14534 2746
rect 14238 2692 14294 2694
rect 14318 2692 14374 2694
rect 14398 2692 14454 2694
rect 14478 2692 14534 2694
rect 19551 13626 19607 13628
rect 19631 13626 19687 13628
rect 19711 13626 19767 13628
rect 19791 13626 19847 13628
rect 19551 13574 19597 13626
rect 19597 13574 19607 13626
rect 19631 13574 19661 13626
rect 19661 13574 19673 13626
rect 19673 13574 19687 13626
rect 19711 13574 19725 13626
rect 19725 13574 19737 13626
rect 19737 13574 19767 13626
rect 19791 13574 19801 13626
rect 19801 13574 19847 13626
rect 19551 13572 19607 13574
rect 19631 13572 19687 13574
rect 19711 13572 19767 13574
rect 19791 13572 19847 13574
rect 21546 17720 21602 17776
rect 21546 17060 21602 17096
rect 21546 17040 21548 17060
rect 21548 17040 21600 17060
rect 21600 17040 21602 17060
rect 20211 14170 20267 14172
rect 20291 14170 20347 14172
rect 20371 14170 20427 14172
rect 20451 14170 20507 14172
rect 20211 14118 20257 14170
rect 20257 14118 20267 14170
rect 20291 14118 20321 14170
rect 20321 14118 20333 14170
rect 20333 14118 20347 14170
rect 20371 14118 20385 14170
rect 20385 14118 20397 14170
rect 20397 14118 20427 14170
rect 20451 14118 20461 14170
rect 20461 14118 20507 14170
rect 20211 14116 20267 14118
rect 20291 14116 20347 14118
rect 20371 14116 20427 14118
rect 20451 14116 20507 14118
rect 20211 13082 20267 13084
rect 20291 13082 20347 13084
rect 20371 13082 20427 13084
rect 20451 13082 20507 13084
rect 20211 13030 20257 13082
rect 20257 13030 20267 13082
rect 20291 13030 20321 13082
rect 20321 13030 20333 13082
rect 20333 13030 20347 13082
rect 20371 13030 20385 13082
rect 20385 13030 20397 13082
rect 20397 13030 20427 13082
rect 20451 13030 20461 13082
rect 20461 13030 20507 13082
rect 20211 13028 20267 13030
rect 20291 13028 20347 13030
rect 20371 13028 20427 13030
rect 20451 13028 20507 13030
rect 22006 19080 22062 19136
rect 22006 18400 22062 18456
rect 22006 16360 22062 16416
rect 22006 15680 22062 15736
rect 22006 15000 22062 15056
rect 22006 14356 22008 14376
rect 22008 14356 22060 14376
rect 22060 14356 22062 14376
rect 22006 14320 22062 14356
rect 22006 13640 22062 13696
rect 22006 12960 22062 13016
rect 19551 12538 19607 12540
rect 19631 12538 19687 12540
rect 19711 12538 19767 12540
rect 19791 12538 19847 12540
rect 19551 12486 19597 12538
rect 19597 12486 19607 12538
rect 19631 12486 19661 12538
rect 19661 12486 19673 12538
rect 19673 12486 19687 12538
rect 19711 12486 19725 12538
rect 19725 12486 19737 12538
rect 19737 12486 19767 12538
rect 19791 12486 19801 12538
rect 19801 12486 19847 12538
rect 19551 12484 19607 12486
rect 19631 12484 19687 12486
rect 19711 12484 19767 12486
rect 19791 12484 19847 12486
rect 20211 11994 20267 11996
rect 20291 11994 20347 11996
rect 20371 11994 20427 11996
rect 20451 11994 20507 11996
rect 20211 11942 20257 11994
rect 20257 11942 20267 11994
rect 20291 11942 20321 11994
rect 20321 11942 20333 11994
rect 20333 11942 20347 11994
rect 20371 11942 20385 11994
rect 20385 11942 20397 11994
rect 20397 11942 20427 11994
rect 20451 11942 20461 11994
rect 20461 11942 20507 11994
rect 20211 11940 20267 11942
rect 20291 11940 20347 11942
rect 20371 11940 20427 11942
rect 20451 11940 20507 11942
rect 19551 11450 19607 11452
rect 19631 11450 19687 11452
rect 19711 11450 19767 11452
rect 19791 11450 19847 11452
rect 19551 11398 19597 11450
rect 19597 11398 19607 11450
rect 19631 11398 19661 11450
rect 19661 11398 19673 11450
rect 19673 11398 19687 11450
rect 19711 11398 19725 11450
rect 19725 11398 19737 11450
rect 19737 11398 19767 11450
rect 19791 11398 19801 11450
rect 19801 11398 19847 11450
rect 19551 11396 19607 11398
rect 19631 11396 19687 11398
rect 19711 11396 19767 11398
rect 19791 11396 19847 11398
rect 20211 10906 20267 10908
rect 20291 10906 20347 10908
rect 20371 10906 20427 10908
rect 20451 10906 20507 10908
rect 20211 10854 20257 10906
rect 20257 10854 20267 10906
rect 20291 10854 20321 10906
rect 20321 10854 20333 10906
rect 20333 10854 20347 10906
rect 20371 10854 20385 10906
rect 20385 10854 20397 10906
rect 20397 10854 20427 10906
rect 20451 10854 20461 10906
rect 20461 10854 20507 10906
rect 20211 10852 20267 10854
rect 20291 10852 20347 10854
rect 20371 10852 20427 10854
rect 20451 10852 20507 10854
rect 19551 10362 19607 10364
rect 19631 10362 19687 10364
rect 19711 10362 19767 10364
rect 19791 10362 19847 10364
rect 19551 10310 19597 10362
rect 19597 10310 19607 10362
rect 19631 10310 19661 10362
rect 19661 10310 19673 10362
rect 19673 10310 19687 10362
rect 19711 10310 19725 10362
rect 19725 10310 19737 10362
rect 19737 10310 19767 10362
rect 19791 10310 19801 10362
rect 19801 10310 19847 10362
rect 19551 10308 19607 10310
rect 19631 10308 19687 10310
rect 19711 10308 19767 10310
rect 19791 10308 19847 10310
rect 22006 12280 22062 12336
rect 22006 11600 22062 11656
rect 22006 10920 22062 10976
rect 22006 10240 22062 10296
rect 20211 9818 20267 9820
rect 20291 9818 20347 9820
rect 20371 9818 20427 9820
rect 20451 9818 20507 9820
rect 20211 9766 20257 9818
rect 20257 9766 20267 9818
rect 20291 9766 20321 9818
rect 20321 9766 20333 9818
rect 20333 9766 20347 9818
rect 20371 9766 20385 9818
rect 20385 9766 20397 9818
rect 20397 9766 20427 9818
rect 20451 9766 20461 9818
rect 20461 9766 20507 9818
rect 20211 9764 20267 9766
rect 20291 9764 20347 9766
rect 20371 9764 20427 9766
rect 20451 9764 20507 9766
rect 19551 9274 19607 9276
rect 19631 9274 19687 9276
rect 19711 9274 19767 9276
rect 19791 9274 19847 9276
rect 19551 9222 19597 9274
rect 19597 9222 19607 9274
rect 19631 9222 19661 9274
rect 19661 9222 19673 9274
rect 19673 9222 19687 9274
rect 19711 9222 19725 9274
rect 19725 9222 19737 9274
rect 19737 9222 19767 9274
rect 19791 9222 19801 9274
rect 19801 9222 19847 9274
rect 19551 9220 19607 9222
rect 19631 9220 19687 9222
rect 19711 9220 19767 9222
rect 19791 9220 19847 9222
rect 20211 8730 20267 8732
rect 20291 8730 20347 8732
rect 20371 8730 20427 8732
rect 20451 8730 20507 8732
rect 20211 8678 20257 8730
rect 20257 8678 20267 8730
rect 20291 8678 20321 8730
rect 20321 8678 20333 8730
rect 20333 8678 20347 8730
rect 20371 8678 20385 8730
rect 20385 8678 20397 8730
rect 20397 8678 20427 8730
rect 20451 8678 20461 8730
rect 20461 8678 20507 8730
rect 20211 8676 20267 8678
rect 20291 8676 20347 8678
rect 20371 8676 20427 8678
rect 20451 8676 20507 8678
rect 19551 8186 19607 8188
rect 19631 8186 19687 8188
rect 19711 8186 19767 8188
rect 19791 8186 19847 8188
rect 19551 8134 19597 8186
rect 19597 8134 19607 8186
rect 19631 8134 19661 8186
rect 19661 8134 19673 8186
rect 19673 8134 19687 8186
rect 19711 8134 19725 8186
rect 19725 8134 19737 8186
rect 19737 8134 19767 8186
rect 19791 8134 19801 8186
rect 19801 8134 19847 8186
rect 19551 8132 19607 8134
rect 19631 8132 19687 8134
rect 19711 8132 19767 8134
rect 19791 8132 19847 8134
rect 19551 7098 19607 7100
rect 19631 7098 19687 7100
rect 19711 7098 19767 7100
rect 19791 7098 19847 7100
rect 19551 7046 19597 7098
rect 19597 7046 19607 7098
rect 19631 7046 19661 7098
rect 19661 7046 19673 7098
rect 19673 7046 19687 7098
rect 19711 7046 19725 7098
rect 19725 7046 19737 7098
rect 19737 7046 19767 7098
rect 19791 7046 19801 7098
rect 19801 7046 19847 7098
rect 19551 7044 19607 7046
rect 19631 7044 19687 7046
rect 19711 7044 19767 7046
rect 19791 7044 19847 7046
rect 20211 7642 20267 7644
rect 20291 7642 20347 7644
rect 20371 7642 20427 7644
rect 20451 7642 20507 7644
rect 20211 7590 20257 7642
rect 20257 7590 20267 7642
rect 20291 7590 20321 7642
rect 20321 7590 20333 7642
rect 20333 7590 20347 7642
rect 20371 7590 20385 7642
rect 20385 7590 20397 7642
rect 20397 7590 20427 7642
rect 20451 7590 20461 7642
rect 20461 7590 20507 7642
rect 20211 7588 20267 7590
rect 20291 7588 20347 7590
rect 20371 7588 20427 7590
rect 20451 7588 20507 7590
rect 19551 6010 19607 6012
rect 19631 6010 19687 6012
rect 19711 6010 19767 6012
rect 19791 6010 19847 6012
rect 19551 5958 19597 6010
rect 19597 5958 19607 6010
rect 19631 5958 19661 6010
rect 19661 5958 19673 6010
rect 19673 5958 19687 6010
rect 19711 5958 19725 6010
rect 19725 5958 19737 6010
rect 19737 5958 19767 6010
rect 19791 5958 19801 6010
rect 19801 5958 19847 6010
rect 19551 5956 19607 5958
rect 19631 5956 19687 5958
rect 19711 5956 19767 5958
rect 19791 5956 19847 5958
rect 19551 4922 19607 4924
rect 19631 4922 19687 4924
rect 19711 4922 19767 4924
rect 19791 4922 19847 4924
rect 19551 4870 19597 4922
rect 19597 4870 19607 4922
rect 19631 4870 19661 4922
rect 19661 4870 19673 4922
rect 19673 4870 19687 4922
rect 19711 4870 19725 4922
rect 19725 4870 19737 4922
rect 19737 4870 19767 4922
rect 19791 4870 19801 4922
rect 19801 4870 19847 4922
rect 19551 4868 19607 4870
rect 19631 4868 19687 4870
rect 19711 4868 19767 4870
rect 19791 4868 19847 4870
rect 20211 6554 20267 6556
rect 20291 6554 20347 6556
rect 20371 6554 20427 6556
rect 20451 6554 20507 6556
rect 20211 6502 20257 6554
rect 20257 6502 20267 6554
rect 20291 6502 20321 6554
rect 20321 6502 20333 6554
rect 20333 6502 20347 6554
rect 20371 6502 20385 6554
rect 20385 6502 20397 6554
rect 20397 6502 20427 6554
rect 20451 6502 20461 6554
rect 20461 6502 20507 6554
rect 20211 6500 20267 6502
rect 20291 6500 20347 6502
rect 20371 6500 20427 6502
rect 20451 6500 20507 6502
rect 20211 5466 20267 5468
rect 20291 5466 20347 5468
rect 20371 5466 20427 5468
rect 20451 5466 20507 5468
rect 20211 5414 20257 5466
rect 20257 5414 20267 5466
rect 20291 5414 20321 5466
rect 20321 5414 20333 5466
rect 20333 5414 20347 5466
rect 20371 5414 20385 5466
rect 20385 5414 20397 5466
rect 20397 5414 20427 5466
rect 20451 5414 20461 5466
rect 20461 5414 20507 5466
rect 20211 5412 20267 5414
rect 20291 5412 20347 5414
rect 20371 5412 20427 5414
rect 20451 5412 20507 5414
rect 21914 9560 21970 9616
rect 21914 8880 21970 8936
rect 21546 8200 21602 8256
rect 21914 7520 21970 7576
rect 22006 6840 22062 6896
rect 21546 6180 21602 6216
rect 21546 6160 21548 6180
rect 21548 6160 21600 6180
rect 21600 6160 21602 6180
rect 22006 5480 22062 5536
rect 22006 4800 22062 4856
rect 20211 4378 20267 4380
rect 20291 4378 20347 4380
rect 20371 4378 20427 4380
rect 20451 4378 20507 4380
rect 20211 4326 20257 4378
rect 20257 4326 20267 4378
rect 20291 4326 20321 4378
rect 20321 4326 20333 4378
rect 20333 4326 20347 4378
rect 20371 4326 20385 4378
rect 20385 4326 20397 4378
rect 20397 4326 20427 4378
rect 20451 4326 20461 4378
rect 20461 4326 20507 4378
rect 20211 4324 20267 4326
rect 20291 4324 20347 4326
rect 20371 4324 20427 4326
rect 20451 4324 20507 4326
rect 19551 3834 19607 3836
rect 19631 3834 19687 3836
rect 19711 3834 19767 3836
rect 19791 3834 19847 3836
rect 19551 3782 19597 3834
rect 19597 3782 19607 3834
rect 19631 3782 19661 3834
rect 19661 3782 19673 3834
rect 19673 3782 19687 3834
rect 19711 3782 19725 3834
rect 19725 3782 19737 3834
rect 19737 3782 19767 3834
rect 19791 3782 19801 3834
rect 19801 3782 19847 3834
rect 19551 3780 19607 3782
rect 19631 3780 19687 3782
rect 19711 3780 19767 3782
rect 19791 3780 19847 3782
rect 20211 3290 20267 3292
rect 20291 3290 20347 3292
rect 20371 3290 20427 3292
rect 20451 3290 20507 3292
rect 20211 3238 20257 3290
rect 20257 3238 20267 3290
rect 20291 3238 20321 3290
rect 20321 3238 20333 3290
rect 20333 3238 20347 3290
rect 20371 3238 20385 3290
rect 20385 3238 20397 3290
rect 20397 3238 20427 3290
rect 20451 3238 20461 3290
rect 20461 3238 20507 3290
rect 20211 3236 20267 3238
rect 20291 3236 20347 3238
rect 20371 3236 20427 3238
rect 20451 3236 20507 3238
rect 19551 2746 19607 2748
rect 19631 2746 19687 2748
rect 19711 2746 19767 2748
rect 19791 2746 19847 2748
rect 19551 2694 19597 2746
rect 19597 2694 19607 2746
rect 19631 2694 19661 2746
rect 19661 2694 19673 2746
rect 19673 2694 19687 2746
rect 19711 2694 19725 2746
rect 19725 2694 19737 2746
rect 19737 2694 19767 2746
rect 19791 2694 19801 2746
rect 19801 2694 19847 2746
rect 19551 2692 19607 2694
rect 19631 2692 19687 2694
rect 19711 2692 19767 2694
rect 19791 2692 19847 2694
rect 22006 4120 22062 4176
rect 14898 2202 14954 2204
rect 14978 2202 15034 2204
rect 15058 2202 15114 2204
rect 15138 2202 15194 2204
rect 14898 2150 14944 2202
rect 14944 2150 14954 2202
rect 14978 2150 15008 2202
rect 15008 2150 15020 2202
rect 15020 2150 15034 2202
rect 15058 2150 15072 2202
rect 15072 2150 15084 2202
rect 15084 2150 15114 2202
rect 15138 2150 15148 2202
rect 15148 2150 15194 2202
rect 14898 2148 14954 2150
rect 14978 2148 15034 2150
rect 15058 2148 15114 2150
rect 15138 2148 15194 2150
rect 20211 2202 20267 2204
rect 20291 2202 20347 2204
rect 20371 2202 20427 2204
rect 20451 2202 20507 2204
rect 20211 2150 20257 2202
rect 20257 2150 20267 2202
rect 20291 2150 20321 2202
rect 20321 2150 20333 2202
rect 20333 2150 20347 2202
rect 20371 2150 20385 2202
rect 20385 2150 20397 2202
rect 20397 2150 20427 2202
rect 20451 2150 20461 2202
rect 20461 2150 20507 2202
rect 20211 2148 20267 2150
rect 20291 2148 20347 2150
rect 20371 2148 20427 2150
rect 20451 2148 20507 2150
<< metal3 >>
rect 3602 23424 3918 23425
rect 3602 23360 3608 23424
rect 3672 23360 3688 23424
rect 3752 23360 3768 23424
rect 3832 23360 3848 23424
rect 3912 23360 3918 23424
rect 3602 23359 3918 23360
rect 8915 23424 9231 23425
rect 8915 23360 8921 23424
rect 8985 23360 9001 23424
rect 9065 23360 9081 23424
rect 9145 23360 9161 23424
rect 9225 23360 9231 23424
rect 8915 23359 9231 23360
rect 14228 23424 14544 23425
rect 14228 23360 14234 23424
rect 14298 23360 14314 23424
rect 14378 23360 14394 23424
rect 14458 23360 14474 23424
rect 14538 23360 14544 23424
rect 14228 23359 14544 23360
rect 19541 23424 19857 23425
rect 19541 23360 19547 23424
rect 19611 23360 19627 23424
rect 19691 23360 19707 23424
rect 19771 23360 19787 23424
rect 19851 23360 19857 23424
rect 19541 23359 19857 23360
rect 4262 22880 4578 22881
rect 4262 22816 4268 22880
rect 4332 22816 4348 22880
rect 4412 22816 4428 22880
rect 4492 22816 4508 22880
rect 4572 22816 4578 22880
rect 4262 22815 4578 22816
rect 9575 22880 9891 22881
rect 9575 22816 9581 22880
rect 9645 22816 9661 22880
rect 9725 22816 9741 22880
rect 9805 22816 9821 22880
rect 9885 22816 9891 22880
rect 9575 22815 9891 22816
rect 14888 22880 15204 22881
rect 14888 22816 14894 22880
rect 14958 22816 14974 22880
rect 15038 22816 15054 22880
rect 15118 22816 15134 22880
rect 15198 22816 15204 22880
rect 14888 22815 15204 22816
rect 20201 22880 20517 22881
rect 20201 22816 20207 22880
rect 20271 22816 20287 22880
rect 20351 22816 20367 22880
rect 20431 22816 20447 22880
rect 20511 22816 20517 22880
rect 20201 22815 20517 22816
rect 841 22674 907 22677
rect 798 22672 907 22674
rect 798 22616 846 22672
rect 902 22616 907 22672
rect 798 22611 907 22616
rect 798 22568 858 22611
rect 0 22478 858 22568
rect 0 22448 800 22478
rect 3602 22336 3918 22337
rect 3602 22272 3608 22336
rect 3672 22272 3688 22336
rect 3752 22272 3768 22336
rect 3832 22272 3848 22336
rect 3912 22272 3918 22336
rect 3602 22271 3918 22272
rect 8915 22336 9231 22337
rect 8915 22272 8921 22336
rect 8985 22272 9001 22336
rect 9065 22272 9081 22336
rect 9145 22272 9161 22336
rect 9225 22272 9231 22336
rect 8915 22271 9231 22272
rect 14228 22336 14544 22337
rect 14228 22272 14234 22336
rect 14298 22272 14314 22336
rect 14378 22272 14394 22336
rect 14458 22272 14474 22336
rect 14538 22272 14544 22336
rect 14228 22271 14544 22272
rect 19541 22336 19857 22337
rect 19541 22272 19547 22336
rect 19611 22272 19627 22336
rect 19691 22272 19707 22336
rect 19771 22272 19787 22336
rect 19851 22272 19857 22336
rect 19541 22271 19857 22272
rect 841 21994 907 21997
rect 798 21992 907 21994
rect 798 21936 846 21992
rect 902 21936 907 21992
rect 798 21931 907 21936
rect 798 21888 858 21931
rect 0 21798 858 21888
rect 0 21768 800 21798
rect 4262 21792 4578 21793
rect 4262 21728 4268 21792
rect 4332 21728 4348 21792
rect 4412 21728 4428 21792
rect 4492 21728 4508 21792
rect 4572 21728 4578 21792
rect 4262 21727 4578 21728
rect 9575 21792 9891 21793
rect 9575 21728 9581 21792
rect 9645 21728 9661 21792
rect 9725 21728 9741 21792
rect 9805 21728 9821 21792
rect 9885 21728 9891 21792
rect 9575 21727 9891 21728
rect 14888 21792 15204 21793
rect 14888 21728 14894 21792
rect 14958 21728 14974 21792
rect 15038 21728 15054 21792
rect 15118 21728 15134 21792
rect 15198 21728 15204 21792
rect 14888 21727 15204 21728
rect 20201 21792 20517 21793
rect 20201 21728 20207 21792
rect 20271 21728 20287 21792
rect 20351 21728 20367 21792
rect 20431 21728 20447 21792
rect 20511 21728 20517 21792
rect 20201 21727 20517 21728
rect 841 21314 907 21317
rect 798 21312 907 21314
rect 798 21256 846 21312
rect 902 21256 907 21312
rect 798 21251 907 21256
rect 798 21208 858 21251
rect 0 21118 858 21208
rect 3602 21248 3918 21249
rect 3602 21184 3608 21248
rect 3672 21184 3688 21248
rect 3752 21184 3768 21248
rect 3832 21184 3848 21248
rect 3912 21184 3918 21248
rect 3602 21183 3918 21184
rect 8915 21248 9231 21249
rect 8915 21184 8921 21248
rect 8985 21184 9001 21248
rect 9065 21184 9081 21248
rect 9145 21184 9161 21248
rect 9225 21184 9231 21248
rect 8915 21183 9231 21184
rect 14228 21248 14544 21249
rect 14228 21184 14234 21248
rect 14298 21184 14314 21248
rect 14378 21184 14394 21248
rect 14458 21184 14474 21248
rect 14538 21184 14544 21248
rect 14228 21183 14544 21184
rect 19541 21248 19857 21249
rect 19541 21184 19547 21248
rect 19611 21184 19627 21248
rect 19691 21184 19707 21248
rect 19771 21184 19787 21248
rect 19851 21184 19857 21248
rect 19541 21183 19857 21184
rect 0 21088 800 21118
rect 4262 20704 4578 20705
rect 4262 20640 4268 20704
rect 4332 20640 4348 20704
rect 4412 20640 4428 20704
rect 4492 20640 4508 20704
rect 4572 20640 4578 20704
rect 4262 20639 4578 20640
rect 9575 20704 9891 20705
rect 9575 20640 9581 20704
rect 9645 20640 9661 20704
rect 9725 20640 9741 20704
rect 9805 20640 9821 20704
rect 9885 20640 9891 20704
rect 9575 20639 9891 20640
rect 14888 20704 15204 20705
rect 14888 20640 14894 20704
rect 14958 20640 14974 20704
rect 15038 20640 15054 20704
rect 15118 20640 15134 20704
rect 15198 20640 15204 20704
rect 14888 20639 15204 20640
rect 20201 20704 20517 20705
rect 20201 20640 20207 20704
rect 20271 20640 20287 20704
rect 20351 20640 20367 20704
rect 20431 20640 20447 20704
rect 20511 20640 20517 20704
rect 20201 20639 20517 20640
rect 0 20498 800 20528
rect 1485 20498 1551 20501
rect 0 20496 1551 20498
rect 0 20440 1490 20496
rect 1546 20440 1551 20496
rect 0 20438 1551 20440
rect 0 20408 800 20438
rect 1485 20435 1551 20438
rect 22001 20498 22067 20501
rect 22668 20498 23468 20528
rect 22001 20496 23468 20498
rect 22001 20440 22006 20496
rect 22062 20440 23468 20496
rect 22001 20438 23468 20440
rect 22001 20435 22067 20438
rect 22668 20408 23468 20438
rect 3602 20160 3918 20161
rect 3602 20096 3608 20160
rect 3672 20096 3688 20160
rect 3752 20096 3768 20160
rect 3832 20096 3848 20160
rect 3912 20096 3918 20160
rect 3602 20095 3918 20096
rect 8915 20160 9231 20161
rect 8915 20096 8921 20160
rect 8985 20096 9001 20160
rect 9065 20096 9081 20160
rect 9145 20096 9161 20160
rect 9225 20096 9231 20160
rect 8915 20095 9231 20096
rect 14228 20160 14544 20161
rect 14228 20096 14234 20160
rect 14298 20096 14314 20160
rect 14378 20096 14394 20160
rect 14458 20096 14474 20160
rect 14538 20096 14544 20160
rect 14228 20095 14544 20096
rect 19541 20160 19857 20161
rect 19541 20096 19547 20160
rect 19611 20096 19627 20160
rect 19691 20096 19707 20160
rect 19771 20096 19787 20160
rect 19851 20096 19857 20160
rect 19541 20095 19857 20096
rect 0 19818 800 19848
rect 22001 19818 22067 19821
rect 22668 19818 23468 19848
rect 0 19728 858 19818
rect 22001 19816 23468 19818
rect 22001 19760 22006 19816
rect 22062 19760 23468 19816
rect 22001 19758 23468 19760
rect 22001 19755 22067 19758
rect 22668 19728 23468 19758
rect 798 19685 858 19728
rect 798 19680 907 19685
rect 798 19624 846 19680
rect 902 19624 907 19680
rect 798 19622 907 19624
rect 841 19619 907 19622
rect 4262 19616 4578 19617
rect 4262 19552 4268 19616
rect 4332 19552 4348 19616
rect 4412 19552 4428 19616
rect 4492 19552 4508 19616
rect 4572 19552 4578 19616
rect 4262 19551 4578 19552
rect 9575 19616 9891 19617
rect 9575 19552 9581 19616
rect 9645 19552 9661 19616
rect 9725 19552 9741 19616
rect 9805 19552 9821 19616
rect 9885 19552 9891 19616
rect 9575 19551 9891 19552
rect 14888 19616 15204 19617
rect 14888 19552 14894 19616
rect 14958 19552 14974 19616
rect 15038 19552 15054 19616
rect 15118 19552 15134 19616
rect 15198 19552 15204 19616
rect 14888 19551 15204 19552
rect 20201 19616 20517 19617
rect 20201 19552 20207 19616
rect 20271 19552 20287 19616
rect 20351 19552 20367 19616
rect 20431 19552 20447 19616
rect 20511 19552 20517 19616
rect 20201 19551 20517 19552
rect 0 19138 800 19168
rect 1485 19138 1551 19141
rect 0 19136 1551 19138
rect 0 19080 1490 19136
rect 1546 19080 1551 19136
rect 0 19078 1551 19080
rect 0 19048 800 19078
rect 1485 19075 1551 19078
rect 22001 19138 22067 19141
rect 22668 19138 23468 19168
rect 22001 19136 23468 19138
rect 22001 19080 22006 19136
rect 22062 19080 23468 19136
rect 22001 19078 23468 19080
rect 22001 19075 22067 19078
rect 3602 19072 3918 19073
rect 3602 19008 3608 19072
rect 3672 19008 3688 19072
rect 3752 19008 3768 19072
rect 3832 19008 3848 19072
rect 3912 19008 3918 19072
rect 3602 19007 3918 19008
rect 8915 19072 9231 19073
rect 8915 19008 8921 19072
rect 8985 19008 9001 19072
rect 9065 19008 9081 19072
rect 9145 19008 9161 19072
rect 9225 19008 9231 19072
rect 8915 19007 9231 19008
rect 14228 19072 14544 19073
rect 14228 19008 14234 19072
rect 14298 19008 14314 19072
rect 14378 19008 14394 19072
rect 14458 19008 14474 19072
rect 14538 19008 14544 19072
rect 14228 19007 14544 19008
rect 19541 19072 19857 19073
rect 19541 19008 19547 19072
rect 19611 19008 19627 19072
rect 19691 19008 19707 19072
rect 19771 19008 19787 19072
rect 19851 19008 19857 19072
rect 22668 19048 23468 19078
rect 19541 19007 19857 19008
rect 841 18594 907 18597
rect 798 18592 907 18594
rect 798 18536 846 18592
rect 902 18536 907 18592
rect 798 18531 907 18536
rect 798 18488 858 18531
rect 0 18398 858 18488
rect 4262 18528 4578 18529
rect 4262 18464 4268 18528
rect 4332 18464 4348 18528
rect 4412 18464 4428 18528
rect 4492 18464 4508 18528
rect 4572 18464 4578 18528
rect 4262 18463 4578 18464
rect 9575 18528 9891 18529
rect 9575 18464 9581 18528
rect 9645 18464 9661 18528
rect 9725 18464 9741 18528
rect 9805 18464 9821 18528
rect 9885 18464 9891 18528
rect 9575 18463 9891 18464
rect 14888 18528 15204 18529
rect 14888 18464 14894 18528
rect 14958 18464 14974 18528
rect 15038 18464 15054 18528
rect 15118 18464 15134 18528
rect 15198 18464 15204 18528
rect 14888 18463 15204 18464
rect 20201 18528 20517 18529
rect 20201 18464 20207 18528
rect 20271 18464 20287 18528
rect 20351 18464 20367 18528
rect 20431 18464 20447 18528
rect 20511 18464 20517 18528
rect 20201 18463 20517 18464
rect 22001 18458 22067 18461
rect 22668 18458 23468 18488
rect 22001 18456 23468 18458
rect 22001 18400 22006 18456
rect 22062 18400 23468 18456
rect 22001 18398 23468 18400
rect 0 18368 800 18398
rect 22001 18395 22067 18398
rect 22668 18368 23468 18398
rect 3602 17984 3918 17985
rect 3602 17920 3608 17984
rect 3672 17920 3688 17984
rect 3752 17920 3768 17984
rect 3832 17920 3848 17984
rect 3912 17920 3918 17984
rect 3602 17919 3918 17920
rect 8915 17984 9231 17985
rect 8915 17920 8921 17984
rect 8985 17920 9001 17984
rect 9065 17920 9081 17984
rect 9145 17920 9161 17984
rect 9225 17920 9231 17984
rect 8915 17919 9231 17920
rect 14228 17984 14544 17985
rect 14228 17920 14234 17984
rect 14298 17920 14314 17984
rect 14378 17920 14394 17984
rect 14458 17920 14474 17984
rect 14538 17920 14544 17984
rect 14228 17919 14544 17920
rect 19541 17984 19857 17985
rect 19541 17920 19547 17984
rect 19611 17920 19627 17984
rect 19691 17920 19707 17984
rect 19771 17920 19787 17984
rect 19851 17920 19857 17984
rect 19541 17919 19857 17920
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 21541 17778 21607 17781
rect 22668 17778 23468 17808
rect 21541 17776 23468 17778
rect 21541 17720 21546 17776
rect 21602 17720 23468 17776
rect 21541 17718 23468 17720
rect 21541 17715 21607 17718
rect 22668 17688 23468 17718
rect 4262 17440 4578 17441
rect 4262 17376 4268 17440
rect 4332 17376 4348 17440
rect 4412 17376 4428 17440
rect 4492 17376 4508 17440
rect 4572 17376 4578 17440
rect 4262 17375 4578 17376
rect 9575 17440 9891 17441
rect 9575 17376 9581 17440
rect 9645 17376 9661 17440
rect 9725 17376 9741 17440
rect 9805 17376 9821 17440
rect 9885 17376 9891 17440
rect 9575 17375 9891 17376
rect 14888 17440 15204 17441
rect 14888 17376 14894 17440
rect 14958 17376 14974 17440
rect 15038 17376 15054 17440
rect 15118 17376 15134 17440
rect 15198 17376 15204 17440
rect 14888 17375 15204 17376
rect 20201 17440 20517 17441
rect 20201 17376 20207 17440
rect 20271 17376 20287 17440
rect 20351 17376 20367 17440
rect 20431 17376 20447 17440
rect 20511 17376 20517 17440
rect 20201 17375 20517 17376
rect 0 17098 800 17128
rect 21541 17098 21607 17101
rect 22668 17098 23468 17128
rect 0 17008 858 17098
rect 21541 17096 23468 17098
rect 21541 17040 21546 17096
rect 21602 17040 23468 17096
rect 21541 17038 23468 17040
rect 21541 17035 21607 17038
rect 22668 17008 23468 17038
rect 798 16965 858 17008
rect 798 16960 907 16965
rect 798 16904 846 16960
rect 902 16904 907 16960
rect 798 16902 907 16904
rect 841 16899 907 16902
rect 3602 16896 3918 16897
rect 3602 16832 3608 16896
rect 3672 16832 3688 16896
rect 3752 16832 3768 16896
rect 3832 16832 3848 16896
rect 3912 16832 3918 16896
rect 3602 16831 3918 16832
rect 8915 16896 9231 16897
rect 8915 16832 8921 16896
rect 8985 16832 9001 16896
rect 9065 16832 9081 16896
rect 9145 16832 9161 16896
rect 9225 16832 9231 16896
rect 8915 16831 9231 16832
rect 14228 16896 14544 16897
rect 14228 16832 14234 16896
rect 14298 16832 14314 16896
rect 14378 16832 14394 16896
rect 14458 16832 14474 16896
rect 14538 16832 14544 16896
rect 14228 16831 14544 16832
rect 19541 16896 19857 16897
rect 19541 16832 19547 16896
rect 19611 16832 19627 16896
rect 19691 16832 19707 16896
rect 19771 16832 19787 16896
rect 19851 16832 19857 16896
rect 19541 16831 19857 16832
rect 841 16554 907 16557
rect 798 16552 907 16554
rect 798 16496 846 16552
rect 902 16496 907 16552
rect 798 16491 907 16496
rect 798 16448 858 16491
rect 0 16358 858 16448
rect 22001 16418 22067 16421
rect 22668 16418 23468 16448
rect 22001 16416 23468 16418
rect 22001 16360 22006 16416
rect 22062 16360 23468 16416
rect 22001 16358 23468 16360
rect 0 16328 800 16358
rect 22001 16355 22067 16358
rect 4262 16352 4578 16353
rect 4262 16288 4268 16352
rect 4332 16288 4348 16352
rect 4412 16288 4428 16352
rect 4492 16288 4508 16352
rect 4572 16288 4578 16352
rect 4262 16287 4578 16288
rect 9575 16352 9891 16353
rect 9575 16288 9581 16352
rect 9645 16288 9661 16352
rect 9725 16288 9741 16352
rect 9805 16288 9821 16352
rect 9885 16288 9891 16352
rect 9575 16287 9891 16288
rect 14888 16352 15204 16353
rect 14888 16288 14894 16352
rect 14958 16288 14974 16352
rect 15038 16288 15054 16352
rect 15118 16288 15134 16352
rect 15198 16288 15204 16352
rect 14888 16287 15204 16288
rect 20201 16352 20517 16353
rect 20201 16288 20207 16352
rect 20271 16288 20287 16352
rect 20351 16288 20367 16352
rect 20431 16288 20447 16352
rect 20511 16288 20517 16352
rect 22668 16328 23468 16358
rect 20201 16287 20517 16288
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 3602 15808 3918 15809
rect 3602 15744 3608 15808
rect 3672 15744 3688 15808
rect 3752 15744 3768 15808
rect 3832 15744 3848 15808
rect 3912 15744 3918 15808
rect 3602 15743 3918 15744
rect 8915 15808 9231 15809
rect 8915 15744 8921 15808
rect 8985 15744 9001 15808
rect 9065 15744 9081 15808
rect 9145 15744 9161 15808
rect 9225 15744 9231 15808
rect 8915 15743 9231 15744
rect 14228 15808 14544 15809
rect 14228 15744 14234 15808
rect 14298 15744 14314 15808
rect 14378 15744 14394 15808
rect 14458 15744 14474 15808
rect 14538 15744 14544 15808
rect 14228 15743 14544 15744
rect 19541 15808 19857 15809
rect 19541 15744 19547 15808
rect 19611 15744 19627 15808
rect 19691 15744 19707 15808
rect 19771 15744 19787 15808
rect 19851 15744 19857 15808
rect 19541 15743 19857 15744
rect 22001 15738 22067 15741
rect 22668 15738 23468 15768
rect 22001 15736 23468 15738
rect 22001 15680 22006 15736
rect 22062 15680 23468 15736
rect 22001 15678 23468 15680
rect 0 15648 800 15678
rect 22001 15675 22067 15678
rect 22668 15648 23468 15678
rect 4262 15264 4578 15265
rect 4262 15200 4268 15264
rect 4332 15200 4348 15264
rect 4412 15200 4428 15264
rect 4492 15200 4508 15264
rect 4572 15200 4578 15264
rect 4262 15199 4578 15200
rect 9575 15264 9891 15265
rect 9575 15200 9581 15264
rect 9645 15200 9661 15264
rect 9725 15200 9741 15264
rect 9805 15200 9821 15264
rect 9885 15200 9891 15264
rect 9575 15199 9891 15200
rect 14888 15264 15204 15265
rect 14888 15200 14894 15264
rect 14958 15200 14974 15264
rect 15038 15200 15054 15264
rect 15118 15200 15134 15264
rect 15198 15200 15204 15264
rect 14888 15199 15204 15200
rect 20201 15264 20517 15265
rect 20201 15200 20207 15264
rect 20271 15200 20287 15264
rect 20351 15200 20367 15264
rect 20431 15200 20447 15264
rect 20511 15200 20517 15264
rect 20201 15199 20517 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 22001 15058 22067 15061
rect 22668 15058 23468 15088
rect 22001 15056 23468 15058
rect 22001 15000 22006 15056
rect 22062 15000 23468 15056
rect 22001 14998 23468 15000
rect 22001 14995 22067 14998
rect 22668 14968 23468 14998
rect 3602 14720 3918 14721
rect 3602 14656 3608 14720
rect 3672 14656 3688 14720
rect 3752 14656 3768 14720
rect 3832 14656 3848 14720
rect 3912 14656 3918 14720
rect 3602 14655 3918 14656
rect 8915 14720 9231 14721
rect 8915 14656 8921 14720
rect 8985 14656 9001 14720
rect 9065 14656 9081 14720
rect 9145 14656 9161 14720
rect 9225 14656 9231 14720
rect 8915 14655 9231 14656
rect 14228 14720 14544 14721
rect 14228 14656 14234 14720
rect 14298 14656 14314 14720
rect 14378 14656 14394 14720
rect 14458 14656 14474 14720
rect 14538 14656 14544 14720
rect 14228 14655 14544 14656
rect 19541 14720 19857 14721
rect 19541 14656 19547 14720
rect 19611 14656 19627 14720
rect 19691 14656 19707 14720
rect 19771 14656 19787 14720
rect 19851 14656 19857 14720
rect 19541 14655 19857 14656
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 22001 14378 22067 14381
rect 22668 14378 23468 14408
rect 22001 14376 23468 14378
rect 22001 14320 22006 14376
rect 22062 14320 23468 14376
rect 22001 14318 23468 14320
rect 0 14288 800 14318
rect 22001 14315 22067 14318
rect 22668 14288 23468 14318
rect 4262 14176 4578 14177
rect 4262 14112 4268 14176
rect 4332 14112 4348 14176
rect 4412 14112 4428 14176
rect 4492 14112 4508 14176
rect 4572 14112 4578 14176
rect 4262 14111 4578 14112
rect 9575 14176 9891 14177
rect 9575 14112 9581 14176
rect 9645 14112 9661 14176
rect 9725 14112 9741 14176
rect 9805 14112 9821 14176
rect 9885 14112 9891 14176
rect 9575 14111 9891 14112
rect 14888 14176 15204 14177
rect 14888 14112 14894 14176
rect 14958 14112 14974 14176
rect 15038 14112 15054 14176
rect 15118 14112 15134 14176
rect 15198 14112 15204 14176
rect 14888 14111 15204 14112
rect 20201 14176 20517 14177
rect 20201 14112 20207 14176
rect 20271 14112 20287 14176
rect 20351 14112 20367 14176
rect 20431 14112 20447 14176
rect 20511 14112 20517 14176
rect 20201 14111 20517 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 22001 13698 22067 13701
rect 22668 13698 23468 13728
rect 22001 13696 23468 13698
rect 22001 13640 22006 13696
rect 22062 13640 23468 13696
rect 22001 13638 23468 13640
rect 22001 13635 22067 13638
rect 3602 13632 3918 13633
rect 3602 13568 3608 13632
rect 3672 13568 3688 13632
rect 3752 13568 3768 13632
rect 3832 13568 3848 13632
rect 3912 13568 3918 13632
rect 3602 13567 3918 13568
rect 8915 13632 9231 13633
rect 8915 13568 8921 13632
rect 8985 13568 9001 13632
rect 9065 13568 9081 13632
rect 9145 13568 9161 13632
rect 9225 13568 9231 13632
rect 8915 13567 9231 13568
rect 14228 13632 14544 13633
rect 14228 13568 14234 13632
rect 14298 13568 14314 13632
rect 14378 13568 14394 13632
rect 14458 13568 14474 13632
rect 14538 13568 14544 13632
rect 14228 13567 14544 13568
rect 19541 13632 19857 13633
rect 19541 13568 19547 13632
rect 19611 13568 19627 13632
rect 19691 13568 19707 13632
rect 19771 13568 19787 13632
rect 19851 13568 19857 13632
rect 22668 13608 23468 13638
rect 19541 13567 19857 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 4262 13088 4578 13089
rect 4262 13024 4268 13088
rect 4332 13024 4348 13088
rect 4412 13024 4428 13088
rect 4492 13024 4508 13088
rect 4572 13024 4578 13088
rect 4262 13023 4578 13024
rect 9575 13088 9891 13089
rect 9575 13024 9581 13088
rect 9645 13024 9661 13088
rect 9725 13024 9741 13088
rect 9805 13024 9821 13088
rect 9885 13024 9891 13088
rect 9575 13023 9891 13024
rect 14888 13088 15204 13089
rect 14888 13024 14894 13088
rect 14958 13024 14974 13088
rect 15038 13024 15054 13088
rect 15118 13024 15134 13088
rect 15198 13024 15204 13088
rect 14888 13023 15204 13024
rect 20201 13088 20517 13089
rect 20201 13024 20207 13088
rect 20271 13024 20287 13088
rect 20351 13024 20367 13088
rect 20431 13024 20447 13088
rect 20511 13024 20517 13088
rect 20201 13023 20517 13024
rect 22001 13018 22067 13021
rect 22668 13018 23468 13048
rect 22001 13016 23468 13018
rect 22001 12960 22006 13016
rect 22062 12960 23468 13016
rect 22001 12958 23468 12960
rect 0 12928 800 12958
rect 22001 12955 22067 12958
rect 22668 12928 23468 12958
rect 3602 12544 3918 12545
rect 3602 12480 3608 12544
rect 3672 12480 3688 12544
rect 3752 12480 3768 12544
rect 3832 12480 3848 12544
rect 3912 12480 3918 12544
rect 3602 12479 3918 12480
rect 8915 12544 9231 12545
rect 8915 12480 8921 12544
rect 8985 12480 9001 12544
rect 9065 12480 9081 12544
rect 9145 12480 9161 12544
rect 9225 12480 9231 12544
rect 8915 12479 9231 12480
rect 14228 12544 14544 12545
rect 14228 12480 14234 12544
rect 14298 12480 14314 12544
rect 14378 12480 14394 12544
rect 14458 12480 14474 12544
rect 14538 12480 14544 12544
rect 14228 12479 14544 12480
rect 19541 12544 19857 12545
rect 19541 12480 19547 12544
rect 19611 12480 19627 12544
rect 19691 12480 19707 12544
rect 19771 12480 19787 12544
rect 19851 12480 19857 12544
rect 19541 12479 19857 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 22001 12338 22067 12341
rect 22668 12338 23468 12368
rect 22001 12336 23468 12338
rect 22001 12280 22006 12336
rect 22062 12280 23468 12336
rect 22001 12278 23468 12280
rect 22001 12275 22067 12278
rect 22668 12248 23468 12278
rect 4262 12000 4578 12001
rect 4262 11936 4268 12000
rect 4332 11936 4348 12000
rect 4412 11936 4428 12000
rect 4492 11936 4508 12000
rect 4572 11936 4578 12000
rect 4262 11935 4578 11936
rect 9575 12000 9891 12001
rect 9575 11936 9581 12000
rect 9645 11936 9661 12000
rect 9725 11936 9741 12000
rect 9805 11936 9821 12000
rect 9885 11936 9891 12000
rect 9575 11935 9891 11936
rect 14888 12000 15204 12001
rect 14888 11936 14894 12000
rect 14958 11936 14974 12000
rect 15038 11936 15054 12000
rect 15118 11936 15134 12000
rect 15198 11936 15204 12000
rect 14888 11935 15204 11936
rect 20201 12000 20517 12001
rect 20201 11936 20207 12000
rect 20271 11936 20287 12000
rect 20351 11936 20367 12000
rect 20431 11936 20447 12000
rect 20511 11936 20517 12000
rect 20201 11935 20517 11936
rect 841 11794 907 11797
rect 798 11792 907 11794
rect 798 11736 846 11792
rect 902 11736 907 11792
rect 798 11731 907 11736
rect 798 11688 858 11731
rect 0 11598 858 11688
rect 22001 11658 22067 11661
rect 22668 11658 23468 11688
rect 22001 11656 23468 11658
rect 22001 11600 22006 11656
rect 22062 11600 23468 11656
rect 22001 11598 23468 11600
rect 0 11568 800 11598
rect 22001 11595 22067 11598
rect 22668 11568 23468 11598
rect 3602 11456 3918 11457
rect 3602 11392 3608 11456
rect 3672 11392 3688 11456
rect 3752 11392 3768 11456
rect 3832 11392 3848 11456
rect 3912 11392 3918 11456
rect 3602 11391 3918 11392
rect 8915 11456 9231 11457
rect 8915 11392 8921 11456
rect 8985 11392 9001 11456
rect 9065 11392 9081 11456
rect 9145 11392 9161 11456
rect 9225 11392 9231 11456
rect 8915 11391 9231 11392
rect 14228 11456 14544 11457
rect 14228 11392 14234 11456
rect 14298 11392 14314 11456
rect 14378 11392 14394 11456
rect 14458 11392 14474 11456
rect 14538 11392 14544 11456
rect 14228 11391 14544 11392
rect 19541 11456 19857 11457
rect 19541 11392 19547 11456
rect 19611 11392 19627 11456
rect 19691 11392 19707 11456
rect 19771 11392 19787 11456
rect 19851 11392 19857 11456
rect 19541 11391 19857 11392
rect 0 10978 800 11008
rect 1669 10978 1735 10981
rect 0 10976 1735 10978
rect 0 10920 1674 10976
rect 1730 10920 1735 10976
rect 0 10918 1735 10920
rect 0 10888 800 10918
rect 1669 10915 1735 10918
rect 22001 10978 22067 10981
rect 22668 10978 23468 11008
rect 22001 10976 23468 10978
rect 22001 10920 22006 10976
rect 22062 10920 23468 10976
rect 22001 10918 23468 10920
rect 22001 10915 22067 10918
rect 4262 10912 4578 10913
rect 4262 10848 4268 10912
rect 4332 10848 4348 10912
rect 4412 10848 4428 10912
rect 4492 10848 4508 10912
rect 4572 10848 4578 10912
rect 4262 10847 4578 10848
rect 9575 10912 9891 10913
rect 9575 10848 9581 10912
rect 9645 10848 9661 10912
rect 9725 10848 9741 10912
rect 9805 10848 9821 10912
rect 9885 10848 9891 10912
rect 9575 10847 9891 10848
rect 14888 10912 15204 10913
rect 14888 10848 14894 10912
rect 14958 10848 14974 10912
rect 15038 10848 15054 10912
rect 15118 10848 15134 10912
rect 15198 10848 15204 10912
rect 14888 10847 15204 10848
rect 20201 10912 20517 10913
rect 20201 10848 20207 10912
rect 20271 10848 20287 10912
rect 20351 10848 20367 10912
rect 20431 10848 20447 10912
rect 20511 10848 20517 10912
rect 22668 10888 23468 10918
rect 20201 10847 20517 10848
rect 3602 10368 3918 10369
rect 0 10298 800 10328
rect 3602 10304 3608 10368
rect 3672 10304 3688 10368
rect 3752 10304 3768 10368
rect 3832 10304 3848 10368
rect 3912 10304 3918 10368
rect 3602 10303 3918 10304
rect 8915 10368 9231 10369
rect 8915 10304 8921 10368
rect 8985 10304 9001 10368
rect 9065 10304 9081 10368
rect 9145 10304 9161 10368
rect 9225 10304 9231 10368
rect 8915 10303 9231 10304
rect 14228 10368 14544 10369
rect 14228 10304 14234 10368
rect 14298 10304 14314 10368
rect 14378 10304 14394 10368
rect 14458 10304 14474 10368
rect 14538 10304 14544 10368
rect 14228 10303 14544 10304
rect 19541 10368 19857 10369
rect 19541 10304 19547 10368
rect 19611 10304 19627 10368
rect 19691 10304 19707 10368
rect 19771 10304 19787 10368
rect 19851 10304 19857 10368
rect 19541 10303 19857 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 22001 10298 22067 10301
rect 22668 10298 23468 10328
rect 22001 10296 23468 10298
rect 22001 10240 22006 10296
rect 22062 10240 23468 10296
rect 22001 10238 23468 10240
rect 22001 10235 22067 10238
rect 22668 10208 23468 10238
rect 4262 9824 4578 9825
rect 4262 9760 4268 9824
rect 4332 9760 4348 9824
rect 4412 9760 4428 9824
rect 4492 9760 4508 9824
rect 4572 9760 4578 9824
rect 4262 9759 4578 9760
rect 9575 9824 9891 9825
rect 9575 9760 9581 9824
rect 9645 9760 9661 9824
rect 9725 9760 9741 9824
rect 9805 9760 9821 9824
rect 9885 9760 9891 9824
rect 9575 9759 9891 9760
rect 14888 9824 15204 9825
rect 14888 9760 14894 9824
rect 14958 9760 14974 9824
rect 15038 9760 15054 9824
rect 15118 9760 15134 9824
rect 15198 9760 15204 9824
rect 14888 9759 15204 9760
rect 20201 9824 20517 9825
rect 20201 9760 20207 9824
rect 20271 9760 20287 9824
rect 20351 9760 20367 9824
rect 20431 9760 20447 9824
rect 20511 9760 20517 9824
rect 20201 9759 20517 9760
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 21909 9618 21975 9621
rect 22668 9618 23468 9648
rect 21909 9616 23468 9618
rect 21909 9560 21914 9616
rect 21970 9560 23468 9616
rect 21909 9558 23468 9560
rect 21909 9555 21975 9558
rect 22668 9528 23468 9558
rect 3602 9280 3918 9281
rect 3602 9216 3608 9280
rect 3672 9216 3688 9280
rect 3752 9216 3768 9280
rect 3832 9216 3848 9280
rect 3912 9216 3918 9280
rect 3602 9215 3918 9216
rect 8915 9280 9231 9281
rect 8915 9216 8921 9280
rect 8985 9216 9001 9280
rect 9065 9216 9081 9280
rect 9145 9216 9161 9280
rect 9225 9216 9231 9280
rect 8915 9215 9231 9216
rect 14228 9280 14544 9281
rect 14228 9216 14234 9280
rect 14298 9216 14314 9280
rect 14378 9216 14394 9280
rect 14458 9216 14474 9280
rect 14538 9216 14544 9280
rect 14228 9215 14544 9216
rect 19541 9280 19857 9281
rect 19541 9216 19547 9280
rect 19611 9216 19627 9280
rect 19691 9216 19707 9280
rect 19771 9216 19787 9280
rect 19851 9216 19857 9280
rect 19541 9215 19857 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 21909 8938 21975 8941
rect 22668 8938 23468 8968
rect 21909 8936 23468 8938
rect 21909 8880 21914 8936
rect 21970 8880 23468 8936
rect 21909 8878 23468 8880
rect 0 8848 800 8878
rect 21909 8875 21975 8878
rect 22668 8848 23468 8878
rect 4262 8736 4578 8737
rect 4262 8672 4268 8736
rect 4332 8672 4348 8736
rect 4412 8672 4428 8736
rect 4492 8672 4508 8736
rect 4572 8672 4578 8736
rect 4262 8671 4578 8672
rect 9575 8736 9891 8737
rect 9575 8672 9581 8736
rect 9645 8672 9661 8736
rect 9725 8672 9741 8736
rect 9805 8672 9821 8736
rect 9885 8672 9891 8736
rect 9575 8671 9891 8672
rect 14888 8736 15204 8737
rect 14888 8672 14894 8736
rect 14958 8672 14974 8736
rect 15038 8672 15054 8736
rect 15118 8672 15134 8736
rect 15198 8672 15204 8736
rect 14888 8671 15204 8672
rect 20201 8736 20517 8737
rect 20201 8672 20207 8736
rect 20271 8672 20287 8736
rect 20351 8672 20367 8736
rect 20431 8672 20447 8736
rect 20511 8672 20517 8736
rect 20201 8671 20517 8672
rect 0 8258 800 8288
rect 1485 8258 1551 8261
rect 0 8256 1551 8258
rect 0 8200 1490 8256
rect 1546 8200 1551 8256
rect 0 8198 1551 8200
rect 0 8168 800 8198
rect 1485 8195 1551 8198
rect 21541 8258 21607 8261
rect 22668 8258 23468 8288
rect 21541 8256 23468 8258
rect 21541 8200 21546 8256
rect 21602 8200 23468 8256
rect 21541 8198 23468 8200
rect 21541 8195 21607 8198
rect 3602 8192 3918 8193
rect 3602 8128 3608 8192
rect 3672 8128 3688 8192
rect 3752 8128 3768 8192
rect 3832 8128 3848 8192
rect 3912 8128 3918 8192
rect 3602 8127 3918 8128
rect 8915 8192 9231 8193
rect 8915 8128 8921 8192
rect 8985 8128 9001 8192
rect 9065 8128 9081 8192
rect 9145 8128 9161 8192
rect 9225 8128 9231 8192
rect 8915 8127 9231 8128
rect 14228 8192 14544 8193
rect 14228 8128 14234 8192
rect 14298 8128 14314 8192
rect 14378 8128 14394 8192
rect 14458 8128 14474 8192
rect 14538 8128 14544 8192
rect 14228 8127 14544 8128
rect 19541 8192 19857 8193
rect 19541 8128 19547 8192
rect 19611 8128 19627 8192
rect 19691 8128 19707 8192
rect 19771 8128 19787 8192
rect 19851 8128 19857 8192
rect 22668 8168 23468 8198
rect 19541 8127 19857 8128
rect 4262 7648 4578 7649
rect 0 7578 800 7608
rect 4262 7584 4268 7648
rect 4332 7584 4348 7648
rect 4412 7584 4428 7648
rect 4492 7584 4508 7648
rect 4572 7584 4578 7648
rect 4262 7583 4578 7584
rect 9575 7648 9891 7649
rect 9575 7584 9581 7648
rect 9645 7584 9661 7648
rect 9725 7584 9741 7648
rect 9805 7584 9821 7648
rect 9885 7584 9891 7648
rect 9575 7583 9891 7584
rect 14888 7648 15204 7649
rect 14888 7584 14894 7648
rect 14958 7584 14974 7648
rect 15038 7584 15054 7648
rect 15118 7584 15134 7648
rect 15198 7584 15204 7648
rect 14888 7583 15204 7584
rect 20201 7648 20517 7649
rect 20201 7584 20207 7648
rect 20271 7584 20287 7648
rect 20351 7584 20367 7648
rect 20431 7584 20447 7648
rect 20511 7584 20517 7648
rect 20201 7583 20517 7584
rect 21909 7578 21975 7581
rect 22668 7578 23468 7608
rect 0 7488 858 7578
rect 21909 7576 23468 7578
rect 21909 7520 21914 7576
rect 21970 7520 23468 7576
rect 21909 7518 23468 7520
rect 21909 7515 21975 7518
rect 22668 7488 23468 7518
rect 798 7445 858 7488
rect 798 7440 907 7445
rect 798 7384 846 7440
rect 902 7384 907 7440
rect 798 7382 907 7384
rect 841 7379 907 7382
rect 3602 7104 3918 7105
rect 3602 7040 3608 7104
rect 3672 7040 3688 7104
rect 3752 7040 3768 7104
rect 3832 7040 3848 7104
rect 3912 7040 3918 7104
rect 3602 7039 3918 7040
rect 8915 7104 9231 7105
rect 8915 7040 8921 7104
rect 8985 7040 9001 7104
rect 9065 7040 9081 7104
rect 9145 7040 9161 7104
rect 9225 7040 9231 7104
rect 8915 7039 9231 7040
rect 14228 7104 14544 7105
rect 14228 7040 14234 7104
rect 14298 7040 14314 7104
rect 14378 7040 14394 7104
rect 14458 7040 14474 7104
rect 14538 7040 14544 7104
rect 14228 7039 14544 7040
rect 19541 7104 19857 7105
rect 19541 7040 19547 7104
rect 19611 7040 19627 7104
rect 19691 7040 19707 7104
rect 19771 7040 19787 7104
rect 19851 7040 19857 7104
rect 19541 7039 19857 7040
rect 0 6898 800 6928
rect 1669 6898 1735 6901
rect 0 6896 1735 6898
rect 0 6840 1674 6896
rect 1730 6840 1735 6896
rect 0 6838 1735 6840
rect 0 6808 800 6838
rect 1669 6835 1735 6838
rect 22001 6898 22067 6901
rect 22668 6898 23468 6928
rect 22001 6896 23468 6898
rect 22001 6840 22006 6896
rect 22062 6840 23468 6896
rect 22001 6838 23468 6840
rect 22001 6835 22067 6838
rect 22668 6808 23468 6838
rect 4262 6560 4578 6561
rect 4262 6496 4268 6560
rect 4332 6496 4348 6560
rect 4412 6496 4428 6560
rect 4492 6496 4508 6560
rect 4572 6496 4578 6560
rect 4262 6495 4578 6496
rect 9575 6560 9891 6561
rect 9575 6496 9581 6560
rect 9645 6496 9661 6560
rect 9725 6496 9741 6560
rect 9805 6496 9821 6560
rect 9885 6496 9891 6560
rect 9575 6495 9891 6496
rect 14888 6560 15204 6561
rect 14888 6496 14894 6560
rect 14958 6496 14974 6560
rect 15038 6496 15054 6560
rect 15118 6496 15134 6560
rect 15198 6496 15204 6560
rect 14888 6495 15204 6496
rect 20201 6560 20517 6561
rect 20201 6496 20207 6560
rect 20271 6496 20287 6560
rect 20351 6496 20367 6560
rect 20431 6496 20447 6560
rect 20511 6496 20517 6560
rect 20201 6495 20517 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 21541 6218 21607 6221
rect 22668 6218 23468 6248
rect 21541 6216 23468 6218
rect 21541 6160 21546 6216
rect 21602 6160 23468 6216
rect 21541 6158 23468 6160
rect 0 6128 800 6158
rect 21541 6155 21607 6158
rect 22668 6128 23468 6158
rect 3602 6016 3918 6017
rect 3602 5952 3608 6016
rect 3672 5952 3688 6016
rect 3752 5952 3768 6016
rect 3832 5952 3848 6016
rect 3912 5952 3918 6016
rect 3602 5951 3918 5952
rect 8915 6016 9231 6017
rect 8915 5952 8921 6016
rect 8985 5952 9001 6016
rect 9065 5952 9081 6016
rect 9145 5952 9161 6016
rect 9225 5952 9231 6016
rect 8915 5951 9231 5952
rect 14228 6016 14544 6017
rect 14228 5952 14234 6016
rect 14298 5952 14314 6016
rect 14378 5952 14394 6016
rect 14458 5952 14474 6016
rect 14538 5952 14544 6016
rect 14228 5951 14544 5952
rect 19541 6016 19857 6017
rect 19541 5952 19547 6016
rect 19611 5952 19627 6016
rect 19691 5952 19707 6016
rect 19771 5952 19787 6016
rect 19851 5952 19857 6016
rect 19541 5951 19857 5952
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 22001 5538 22067 5541
rect 22668 5538 23468 5568
rect 22001 5536 23468 5538
rect 22001 5480 22006 5536
rect 22062 5480 23468 5536
rect 22001 5478 23468 5480
rect 22001 5475 22067 5478
rect 4262 5472 4578 5473
rect 4262 5408 4268 5472
rect 4332 5408 4348 5472
rect 4412 5408 4428 5472
rect 4492 5408 4508 5472
rect 4572 5408 4578 5472
rect 4262 5407 4578 5408
rect 9575 5472 9891 5473
rect 9575 5408 9581 5472
rect 9645 5408 9661 5472
rect 9725 5408 9741 5472
rect 9805 5408 9821 5472
rect 9885 5408 9891 5472
rect 9575 5407 9891 5408
rect 14888 5472 15204 5473
rect 14888 5408 14894 5472
rect 14958 5408 14974 5472
rect 15038 5408 15054 5472
rect 15118 5408 15134 5472
rect 15198 5408 15204 5472
rect 14888 5407 15204 5408
rect 20201 5472 20517 5473
rect 20201 5408 20207 5472
rect 20271 5408 20287 5472
rect 20351 5408 20367 5472
rect 20431 5408 20447 5472
rect 20511 5408 20517 5472
rect 22668 5448 23468 5478
rect 20201 5407 20517 5408
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 3602 4928 3918 4929
rect 3602 4864 3608 4928
rect 3672 4864 3688 4928
rect 3752 4864 3768 4928
rect 3832 4864 3848 4928
rect 3912 4864 3918 4928
rect 3602 4863 3918 4864
rect 8915 4928 9231 4929
rect 8915 4864 8921 4928
rect 8985 4864 9001 4928
rect 9065 4864 9081 4928
rect 9145 4864 9161 4928
rect 9225 4864 9231 4928
rect 8915 4863 9231 4864
rect 14228 4928 14544 4929
rect 14228 4864 14234 4928
rect 14298 4864 14314 4928
rect 14378 4864 14394 4928
rect 14458 4864 14474 4928
rect 14538 4864 14544 4928
rect 14228 4863 14544 4864
rect 19541 4928 19857 4929
rect 19541 4864 19547 4928
rect 19611 4864 19627 4928
rect 19691 4864 19707 4928
rect 19771 4864 19787 4928
rect 19851 4864 19857 4928
rect 19541 4863 19857 4864
rect 22001 4858 22067 4861
rect 22668 4858 23468 4888
rect 22001 4856 23468 4858
rect 22001 4800 22006 4856
rect 22062 4800 23468 4856
rect 22001 4798 23468 4800
rect 0 4768 800 4798
rect 22001 4795 22067 4798
rect 22668 4768 23468 4798
rect 4262 4384 4578 4385
rect 4262 4320 4268 4384
rect 4332 4320 4348 4384
rect 4412 4320 4428 4384
rect 4492 4320 4508 4384
rect 4572 4320 4578 4384
rect 4262 4319 4578 4320
rect 9575 4384 9891 4385
rect 9575 4320 9581 4384
rect 9645 4320 9661 4384
rect 9725 4320 9741 4384
rect 9805 4320 9821 4384
rect 9885 4320 9891 4384
rect 9575 4319 9891 4320
rect 14888 4384 15204 4385
rect 14888 4320 14894 4384
rect 14958 4320 14974 4384
rect 15038 4320 15054 4384
rect 15118 4320 15134 4384
rect 15198 4320 15204 4384
rect 14888 4319 15204 4320
rect 20201 4384 20517 4385
rect 20201 4320 20207 4384
rect 20271 4320 20287 4384
rect 20351 4320 20367 4384
rect 20431 4320 20447 4384
rect 20511 4320 20517 4384
rect 20201 4319 20517 4320
rect 841 4314 907 4317
rect 798 4312 907 4314
rect 798 4256 846 4312
rect 902 4256 907 4312
rect 798 4251 907 4256
rect 798 4208 858 4251
rect 0 4118 858 4208
rect 22001 4178 22067 4181
rect 22668 4178 23468 4208
rect 22001 4176 23468 4178
rect 22001 4120 22006 4176
rect 22062 4120 23468 4176
rect 22001 4118 23468 4120
rect 0 4088 800 4118
rect 22001 4115 22067 4118
rect 22668 4088 23468 4118
rect 3602 3840 3918 3841
rect 3602 3776 3608 3840
rect 3672 3776 3688 3840
rect 3752 3776 3768 3840
rect 3832 3776 3848 3840
rect 3912 3776 3918 3840
rect 3602 3775 3918 3776
rect 8915 3840 9231 3841
rect 8915 3776 8921 3840
rect 8985 3776 9001 3840
rect 9065 3776 9081 3840
rect 9145 3776 9161 3840
rect 9225 3776 9231 3840
rect 8915 3775 9231 3776
rect 14228 3840 14544 3841
rect 14228 3776 14234 3840
rect 14298 3776 14314 3840
rect 14378 3776 14394 3840
rect 14458 3776 14474 3840
rect 14538 3776 14544 3840
rect 14228 3775 14544 3776
rect 19541 3840 19857 3841
rect 19541 3776 19547 3840
rect 19611 3776 19627 3840
rect 19691 3776 19707 3840
rect 19771 3776 19787 3840
rect 19851 3776 19857 3840
rect 19541 3775 19857 3776
rect 0 3498 800 3528
rect 0 3408 858 3498
rect 798 3365 858 3408
rect 798 3360 907 3365
rect 798 3304 846 3360
rect 902 3304 907 3360
rect 798 3302 907 3304
rect 841 3299 907 3302
rect 4262 3296 4578 3297
rect 4262 3232 4268 3296
rect 4332 3232 4348 3296
rect 4412 3232 4428 3296
rect 4492 3232 4508 3296
rect 4572 3232 4578 3296
rect 4262 3231 4578 3232
rect 9575 3296 9891 3297
rect 9575 3232 9581 3296
rect 9645 3232 9661 3296
rect 9725 3232 9741 3296
rect 9805 3232 9821 3296
rect 9885 3232 9891 3296
rect 9575 3231 9891 3232
rect 14888 3296 15204 3297
rect 14888 3232 14894 3296
rect 14958 3232 14974 3296
rect 15038 3232 15054 3296
rect 15118 3232 15134 3296
rect 15198 3232 15204 3296
rect 14888 3231 15204 3232
rect 20201 3296 20517 3297
rect 20201 3232 20207 3296
rect 20271 3232 20287 3296
rect 20351 3232 20367 3296
rect 20431 3232 20447 3296
rect 20511 3232 20517 3296
rect 20201 3231 20517 3232
rect 3602 2752 3918 2753
rect 3602 2688 3608 2752
rect 3672 2688 3688 2752
rect 3752 2688 3768 2752
rect 3832 2688 3848 2752
rect 3912 2688 3918 2752
rect 3602 2687 3918 2688
rect 8915 2752 9231 2753
rect 8915 2688 8921 2752
rect 8985 2688 9001 2752
rect 9065 2688 9081 2752
rect 9145 2688 9161 2752
rect 9225 2688 9231 2752
rect 8915 2687 9231 2688
rect 14228 2752 14544 2753
rect 14228 2688 14234 2752
rect 14298 2688 14314 2752
rect 14378 2688 14394 2752
rect 14458 2688 14474 2752
rect 14538 2688 14544 2752
rect 14228 2687 14544 2688
rect 19541 2752 19857 2753
rect 19541 2688 19547 2752
rect 19611 2688 19627 2752
rect 19691 2688 19707 2752
rect 19771 2688 19787 2752
rect 19851 2688 19857 2752
rect 19541 2687 19857 2688
rect 4262 2208 4578 2209
rect 4262 2144 4268 2208
rect 4332 2144 4348 2208
rect 4412 2144 4428 2208
rect 4492 2144 4508 2208
rect 4572 2144 4578 2208
rect 4262 2143 4578 2144
rect 9575 2208 9891 2209
rect 9575 2144 9581 2208
rect 9645 2144 9661 2208
rect 9725 2144 9741 2208
rect 9805 2144 9821 2208
rect 9885 2144 9891 2208
rect 9575 2143 9891 2144
rect 14888 2208 15204 2209
rect 14888 2144 14894 2208
rect 14958 2144 14974 2208
rect 15038 2144 15054 2208
rect 15118 2144 15134 2208
rect 15198 2144 15204 2208
rect 14888 2143 15204 2144
rect 20201 2208 20517 2209
rect 20201 2144 20207 2208
rect 20271 2144 20287 2208
rect 20351 2144 20367 2208
rect 20431 2144 20447 2208
rect 20511 2144 20517 2208
rect 20201 2143 20517 2144
<< via3 >>
rect 3608 23420 3672 23424
rect 3608 23364 3612 23420
rect 3612 23364 3668 23420
rect 3668 23364 3672 23420
rect 3608 23360 3672 23364
rect 3688 23420 3752 23424
rect 3688 23364 3692 23420
rect 3692 23364 3748 23420
rect 3748 23364 3752 23420
rect 3688 23360 3752 23364
rect 3768 23420 3832 23424
rect 3768 23364 3772 23420
rect 3772 23364 3828 23420
rect 3828 23364 3832 23420
rect 3768 23360 3832 23364
rect 3848 23420 3912 23424
rect 3848 23364 3852 23420
rect 3852 23364 3908 23420
rect 3908 23364 3912 23420
rect 3848 23360 3912 23364
rect 8921 23420 8985 23424
rect 8921 23364 8925 23420
rect 8925 23364 8981 23420
rect 8981 23364 8985 23420
rect 8921 23360 8985 23364
rect 9001 23420 9065 23424
rect 9001 23364 9005 23420
rect 9005 23364 9061 23420
rect 9061 23364 9065 23420
rect 9001 23360 9065 23364
rect 9081 23420 9145 23424
rect 9081 23364 9085 23420
rect 9085 23364 9141 23420
rect 9141 23364 9145 23420
rect 9081 23360 9145 23364
rect 9161 23420 9225 23424
rect 9161 23364 9165 23420
rect 9165 23364 9221 23420
rect 9221 23364 9225 23420
rect 9161 23360 9225 23364
rect 14234 23420 14298 23424
rect 14234 23364 14238 23420
rect 14238 23364 14294 23420
rect 14294 23364 14298 23420
rect 14234 23360 14298 23364
rect 14314 23420 14378 23424
rect 14314 23364 14318 23420
rect 14318 23364 14374 23420
rect 14374 23364 14378 23420
rect 14314 23360 14378 23364
rect 14394 23420 14458 23424
rect 14394 23364 14398 23420
rect 14398 23364 14454 23420
rect 14454 23364 14458 23420
rect 14394 23360 14458 23364
rect 14474 23420 14538 23424
rect 14474 23364 14478 23420
rect 14478 23364 14534 23420
rect 14534 23364 14538 23420
rect 14474 23360 14538 23364
rect 19547 23420 19611 23424
rect 19547 23364 19551 23420
rect 19551 23364 19607 23420
rect 19607 23364 19611 23420
rect 19547 23360 19611 23364
rect 19627 23420 19691 23424
rect 19627 23364 19631 23420
rect 19631 23364 19687 23420
rect 19687 23364 19691 23420
rect 19627 23360 19691 23364
rect 19707 23420 19771 23424
rect 19707 23364 19711 23420
rect 19711 23364 19767 23420
rect 19767 23364 19771 23420
rect 19707 23360 19771 23364
rect 19787 23420 19851 23424
rect 19787 23364 19791 23420
rect 19791 23364 19847 23420
rect 19847 23364 19851 23420
rect 19787 23360 19851 23364
rect 4268 22876 4332 22880
rect 4268 22820 4272 22876
rect 4272 22820 4328 22876
rect 4328 22820 4332 22876
rect 4268 22816 4332 22820
rect 4348 22876 4412 22880
rect 4348 22820 4352 22876
rect 4352 22820 4408 22876
rect 4408 22820 4412 22876
rect 4348 22816 4412 22820
rect 4428 22876 4492 22880
rect 4428 22820 4432 22876
rect 4432 22820 4488 22876
rect 4488 22820 4492 22876
rect 4428 22816 4492 22820
rect 4508 22876 4572 22880
rect 4508 22820 4512 22876
rect 4512 22820 4568 22876
rect 4568 22820 4572 22876
rect 4508 22816 4572 22820
rect 9581 22876 9645 22880
rect 9581 22820 9585 22876
rect 9585 22820 9641 22876
rect 9641 22820 9645 22876
rect 9581 22816 9645 22820
rect 9661 22876 9725 22880
rect 9661 22820 9665 22876
rect 9665 22820 9721 22876
rect 9721 22820 9725 22876
rect 9661 22816 9725 22820
rect 9741 22876 9805 22880
rect 9741 22820 9745 22876
rect 9745 22820 9801 22876
rect 9801 22820 9805 22876
rect 9741 22816 9805 22820
rect 9821 22876 9885 22880
rect 9821 22820 9825 22876
rect 9825 22820 9881 22876
rect 9881 22820 9885 22876
rect 9821 22816 9885 22820
rect 14894 22876 14958 22880
rect 14894 22820 14898 22876
rect 14898 22820 14954 22876
rect 14954 22820 14958 22876
rect 14894 22816 14958 22820
rect 14974 22876 15038 22880
rect 14974 22820 14978 22876
rect 14978 22820 15034 22876
rect 15034 22820 15038 22876
rect 14974 22816 15038 22820
rect 15054 22876 15118 22880
rect 15054 22820 15058 22876
rect 15058 22820 15114 22876
rect 15114 22820 15118 22876
rect 15054 22816 15118 22820
rect 15134 22876 15198 22880
rect 15134 22820 15138 22876
rect 15138 22820 15194 22876
rect 15194 22820 15198 22876
rect 15134 22816 15198 22820
rect 20207 22876 20271 22880
rect 20207 22820 20211 22876
rect 20211 22820 20267 22876
rect 20267 22820 20271 22876
rect 20207 22816 20271 22820
rect 20287 22876 20351 22880
rect 20287 22820 20291 22876
rect 20291 22820 20347 22876
rect 20347 22820 20351 22876
rect 20287 22816 20351 22820
rect 20367 22876 20431 22880
rect 20367 22820 20371 22876
rect 20371 22820 20427 22876
rect 20427 22820 20431 22876
rect 20367 22816 20431 22820
rect 20447 22876 20511 22880
rect 20447 22820 20451 22876
rect 20451 22820 20507 22876
rect 20507 22820 20511 22876
rect 20447 22816 20511 22820
rect 3608 22332 3672 22336
rect 3608 22276 3612 22332
rect 3612 22276 3668 22332
rect 3668 22276 3672 22332
rect 3608 22272 3672 22276
rect 3688 22332 3752 22336
rect 3688 22276 3692 22332
rect 3692 22276 3748 22332
rect 3748 22276 3752 22332
rect 3688 22272 3752 22276
rect 3768 22332 3832 22336
rect 3768 22276 3772 22332
rect 3772 22276 3828 22332
rect 3828 22276 3832 22332
rect 3768 22272 3832 22276
rect 3848 22332 3912 22336
rect 3848 22276 3852 22332
rect 3852 22276 3908 22332
rect 3908 22276 3912 22332
rect 3848 22272 3912 22276
rect 8921 22332 8985 22336
rect 8921 22276 8925 22332
rect 8925 22276 8981 22332
rect 8981 22276 8985 22332
rect 8921 22272 8985 22276
rect 9001 22332 9065 22336
rect 9001 22276 9005 22332
rect 9005 22276 9061 22332
rect 9061 22276 9065 22332
rect 9001 22272 9065 22276
rect 9081 22332 9145 22336
rect 9081 22276 9085 22332
rect 9085 22276 9141 22332
rect 9141 22276 9145 22332
rect 9081 22272 9145 22276
rect 9161 22332 9225 22336
rect 9161 22276 9165 22332
rect 9165 22276 9221 22332
rect 9221 22276 9225 22332
rect 9161 22272 9225 22276
rect 14234 22332 14298 22336
rect 14234 22276 14238 22332
rect 14238 22276 14294 22332
rect 14294 22276 14298 22332
rect 14234 22272 14298 22276
rect 14314 22332 14378 22336
rect 14314 22276 14318 22332
rect 14318 22276 14374 22332
rect 14374 22276 14378 22332
rect 14314 22272 14378 22276
rect 14394 22332 14458 22336
rect 14394 22276 14398 22332
rect 14398 22276 14454 22332
rect 14454 22276 14458 22332
rect 14394 22272 14458 22276
rect 14474 22332 14538 22336
rect 14474 22276 14478 22332
rect 14478 22276 14534 22332
rect 14534 22276 14538 22332
rect 14474 22272 14538 22276
rect 19547 22332 19611 22336
rect 19547 22276 19551 22332
rect 19551 22276 19607 22332
rect 19607 22276 19611 22332
rect 19547 22272 19611 22276
rect 19627 22332 19691 22336
rect 19627 22276 19631 22332
rect 19631 22276 19687 22332
rect 19687 22276 19691 22332
rect 19627 22272 19691 22276
rect 19707 22332 19771 22336
rect 19707 22276 19711 22332
rect 19711 22276 19767 22332
rect 19767 22276 19771 22332
rect 19707 22272 19771 22276
rect 19787 22332 19851 22336
rect 19787 22276 19791 22332
rect 19791 22276 19847 22332
rect 19847 22276 19851 22332
rect 19787 22272 19851 22276
rect 4268 21788 4332 21792
rect 4268 21732 4272 21788
rect 4272 21732 4328 21788
rect 4328 21732 4332 21788
rect 4268 21728 4332 21732
rect 4348 21788 4412 21792
rect 4348 21732 4352 21788
rect 4352 21732 4408 21788
rect 4408 21732 4412 21788
rect 4348 21728 4412 21732
rect 4428 21788 4492 21792
rect 4428 21732 4432 21788
rect 4432 21732 4488 21788
rect 4488 21732 4492 21788
rect 4428 21728 4492 21732
rect 4508 21788 4572 21792
rect 4508 21732 4512 21788
rect 4512 21732 4568 21788
rect 4568 21732 4572 21788
rect 4508 21728 4572 21732
rect 9581 21788 9645 21792
rect 9581 21732 9585 21788
rect 9585 21732 9641 21788
rect 9641 21732 9645 21788
rect 9581 21728 9645 21732
rect 9661 21788 9725 21792
rect 9661 21732 9665 21788
rect 9665 21732 9721 21788
rect 9721 21732 9725 21788
rect 9661 21728 9725 21732
rect 9741 21788 9805 21792
rect 9741 21732 9745 21788
rect 9745 21732 9801 21788
rect 9801 21732 9805 21788
rect 9741 21728 9805 21732
rect 9821 21788 9885 21792
rect 9821 21732 9825 21788
rect 9825 21732 9881 21788
rect 9881 21732 9885 21788
rect 9821 21728 9885 21732
rect 14894 21788 14958 21792
rect 14894 21732 14898 21788
rect 14898 21732 14954 21788
rect 14954 21732 14958 21788
rect 14894 21728 14958 21732
rect 14974 21788 15038 21792
rect 14974 21732 14978 21788
rect 14978 21732 15034 21788
rect 15034 21732 15038 21788
rect 14974 21728 15038 21732
rect 15054 21788 15118 21792
rect 15054 21732 15058 21788
rect 15058 21732 15114 21788
rect 15114 21732 15118 21788
rect 15054 21728 15118 21732
rect 15134 21788 15198 21792
rect 15134 21732 15138 21788
rect 15138 21732 15194 21788
rect 15194 21732 15198 21788
rect 15134 21728 15198 21732
rect 20207 21788 20271 21792
rect 20207 21732 20211 21788
rect 20211 21732 20267 21788
rect 20267 21732 20271 21788
rect 20207 21728 20271 21732
rect 20287 21788 20351 21792
rect 20287 21732 20291 21788
rect 20291 21732 20347 21788
rect 20347 21732 20351 21788
rect 20287 21728 20351 21732
rect 20367 21788 20431 21792
rect 20367 21732 20371 21788
rect 20371 21732 20427 21788
rect 20427 21732 20431 21788
rect 20367 21728 20431 21732
rect 20447 21788 20511 21792
rect 20447 21732 20451 21788
rect 20451 21732 20507 21788
rect 20507 21732 20511 21788
rect 20447 21728 20511 21732
rect 3608 21244 3672 21248
rect 3608 21188 3612 21244
rect 3612 21188 3668 21244
rect 3668 21188 3672 21244
rect 3608 21184 3672 21188
rect 3688 21244 3752 21248
rect 3688 21188 3692 21244
rect 3692 21188 3748 21244
rect 3748 21188 3752 21244
rect 3688 21184 3752 21188
rect 3768 21244 3832 21248
rect 3768 21188 3772 21244
rect 3772 21188 3828 21244
rect 3828 21188 3832 21244
rect 3768 21184 3832 21188
rect 3848 21244 3912 21248
rect 3848 21188 3852 21244
rect 3852 21188 3908 21244
rect 3908 21188 3912 21244
rect 3848 21184 3912 21188
rect 8921 21244 8985 21248
rect 8921 21188 8925 21244
rect 8925 21188 8981 21244
rect 8981 21188 8985 21244
rect 8921 21184 8985 21188
rect 9001 21244 9065 21248
rect 9001 21188 9005 21244
rect 9005 21188 9061 21244
rect 9061 21188 9065 21244
rect 9001 21184 9065 21188
rect 9081 21244 9145 21248
rect 9081 21188 9085 21244
rect 9085 21188 9141 21244
rect 9141 21188 9145 21244
rect 9081 21184 9145 21188
rect 9161 21244 9225 21248
rect 9161 21188 9165 21244
rect 9165 21188 9221 21244
rect 9221 21188 9225 21244
rect 9161 21184 9225 21188
rect 14234 21244 14298 21248
rect 14234 21188 14238 21244
rect 14238 21188 14294 21244
rect 14294 21188 14298 21244
rect 14234 21184 14298 21188
rect 14314 21244 14378 21248
rect 14314 21188 14318 21244
rect 14318 21188 14374 21244
rect 14374 21188 14378 21244
rect 14314 21184 14378 21188
rect 14394 21244 14458 21248
rect 14394 21188 14398 21244
rect 14398 21188 14454 21244
rect 14454 21188 14458 21244
rect 14394 21184 14458 21188
rect 14474 21244 14538 21248
rect 14474 21188 14478 21244
rect 14478 21188 14534 21244
rect 14534 21188 14538 21244
rect 14474 21184 14538 21188
rect 19547 21244 19611 21248
rect 19547 21188 19551 21244
rect 19551 21188 19607 21244
rect 19607 21188 19611 21244
rect 19547 21184 19611 21188
rect 19627 21244 19691 21248
rect 19627 21188 19631 21244
rect 19631 21188 19687 21244
rect 19687 21188 19691 21244
rect 19627 21184 19691 21188
rect 19707 21244 19771 21248
rect 19707 21188 19711 21244
rect 19711 21188 19767 21244
rect 19767 21188 19771 21244
rect 19707 21184 19771 21188
rect 19787 21244 19851 21248
rect 19787 21188 19791 21244
rect 19791 21188 19847 21244
rect 19847 21188 19851 21244
rect 19787 21184 19851 21188
rect 4268 20700 4332 20704
rect 4268 20644 4272 20700
rect 4272 20644 4328 20700
rect 4328 20644 4332 20700
rect 4268 20640 4332 20644
rect 4348 20700 4412 20704
rect 4348 20644 4352 20700
rect 4352 20644 4408 20700
rect 4408 20644 4412 20700
rect 4348 20640 4412 20644
rect 4428 20700 4492 20704
rect 4428 20644 4432 20700
rect 4432 20644 4488 20700
rect 4488 20644 4492 20700
rect 4428 20640 4492 20644
rect 4508 20700 4572 20704
rect 4508 20644 4512 20700
rect 4512 20644 4568 20700
rect 4568 20644 4572 20700
rect 4508 20640 4572 20644
rect 9581 20700 9645 20704
rect 9581 20644 9585 20700
rect 9585 20644 9641 20700
rect 9641 20644 9645 20700
rect 9581 20640 9645 20644
rect 9661 20700 9725 20704
rect 9661 20644 9665 20700
rect 9665 20644 9721 20700
rect 9721 20644 9725 20700
rect 9661 20640 9725 20644
rect 9741 20700 9805 20704
rect 9741 20644 9745 20700
rect 9745 20644 9801 20700
rect 9801 20644 9805 20700
rect 9741 20640 9805 20644
rect 9821 20700 9885 20704
rect 9821 20644 9825 20700
rect 9825 20644 9881 20700
rect 9881 20644 9885 20700
rect 9821 20640 9885 20644
rect 14894 20700 14958 20704
rect 14894 20644 14898 20700
rect 14898 20644 14954 20700
rect 14954 20644 14958 20700
rect 14894 20640 14958 20644
rect 14974 20700 15038 20704
rect 14974 20644 14978 20700
rect 14978 20644 15034 20700
rect 15034 20644 15038 20700
rect 14974 20640 15038 20644
rect 15054 20700 15118 20704
rect 15054 20644 15058 20700
rect 15058 20644 15114 20700
rect 15114 20644 15118 20700
rect 15054 20640 15118 20644
rect 15134 20700 15198 20704
rect 15134 20644 15138 20700
rect 15138 20644 15194 20700
rect 15194 20644 15198 20700
rect 15134 20640 15198 20644
rect 20207 20700 20271 20704
rect 20207 20644 20211 20700
rect 20211 20644 20267 20700
rect 20267 20644 20271 20700
rect 20207 20640 20271 20644
rect 20287 20700 20351 20704
rect 20287 20644 20291 20700
rect 20291 20644 20347 20700
rect 20347 20644 20351 20700
rect 20287 20640 20351 20644
rect 20367 20700 20431 20704
rect 20367 20644 20371 20700
rect 20371 20644 20427 20700
rect 20427 20644 20431 20700
rect 20367 20640 20431 20644
rect 20447 20700 20511 20704
rect 20447 20644 20451 20700
rect 20451 20644 20507 20700
rect 20507 20644 20511 20700
rect 20447 20640 20511 20644
rect 3608 20156 3672 20160
rect 3608 20100 3612 20156
rect 3612 20100 3668 20156
rect 3668 20100 3672 20156
rect 3608 20096 3672 20100
rect 3688 20156 3752 20160
rect 3688 20100 3692 20156
rect 3692 20100 3748 20156
rect 3748 20100 3752 20156
rect 3688 20096 3752 20100
rect 3768 20156 3832 20160
rect 3768 20100 3772 20156
rect 3772 20100 3828 20156
rect 3828 20100 3832 20156
rect 3768 20096 3832 20100
rect 3848 20156 3912 20160
rect 3848 20100 3852 20156
rect 3852 20100 3908 20156
rect 3908 20100 3912 20156
rect 3848 20096 3912 20100
rect 8921 20156 8985 20160
rect 8921 20100 8925 20156
rect 8925 20100 8981 20156
rect 8981 20100 8985 20156
rect 8921 20096 8985 20100
rect 9001 20156 9065 20160
rect 9001 20100 9005 20156
rect 9005 20100 9061 20156
rect 9061 20100 9065 20156
rect 9001 20096 9065 20100
rect 9081 20156 9145 20160
rect 9081 20100 9085 20156
rect 9085 20100 9141 20156
rect 9141 20100 9145 20156
rect 9081 20096 9145 20100
rect 9161 20156 9225 20160
rect 9161 20100 9165 20156
rect 9165 20100 9221 20156
rect 9221 20100 9225 20156
rect 9161 20096 9225 20100
rect 14234 20156 14298 20160
rect 14234 20100 14238 20156
rect 14238 20100 14294 20156
rect 14294 20100 14298 20156
rect 14234 20096 14298 20100
rect 14314 20156 14378 20160
rect 14314 20100 14318 20156
rect 14318 20100 14374 20156
rect 14374 20100 14378 20156
rect 14314 20096 14378 20100
rect 14394 20156 14458 20160
rect 14394 20100 14398 20156
rect 14398 20100 14454 20156
rect 14454 20100 14458 20156
rect 14394 20096 14458 20100
rect 14474 20156 14538 20160
rect 14474 20100 14478 20156
rect 14478 20100 14534 20156
rect 14534 20100 14538 20156
rect 14474 20096 14538 20100
rect 19547 20156 19611 20160
rect 19547 20100 19551 20156
rect 19551 20100 19607 20156
rect 19607 20100 19611 20156
rect 19547 20096 19611 20100
rect 19627 20156 19691 20160
rect 19627 20100 19631 20156
rect 19631 20100 19687 20156
rect 19687 20100 19691 20156
rect 19627 20096 19691 20100
rect 19707 20156 19771 20160
rect 19707 20100 19711 20156
rect 19711 20100 19767 20156
rect 19767 20100 19771 20156
rect 19707 20096 19771 20100
rect 19787 20156 19851 20160
rect 19787 20100 19791 20156
rect 19791 20100 19847 20156
rect 19847 20100 19851 20156
rect 19787 20096 19851 20100
rect 4268 19612 4332 19616
rect 4268 19556 4272 19612
rect 4272 19556 4328 19612
rect 4328 19556 4332 19612
rect 4268 19552 4332 19556
rect 4348 19612 4412 19616
rect 4348 19556 4352 19612
rect 4352 19556 4408 19612
rect 4408 19556 4412 19612
rect 4348 19552 4412 19556
rect 4428 19612 4492 19616
rect 4428 19556 4432 19612
rect 4432 19556 4488 19612
rect 4488 19556 4492 19612
rect 4428 19552 4492 19556
rect 4508 19612 4572 19616
rect 4508 19556 4512 19612
rect 4512 19556 4568 19612
rect 4568 19556 4572 19612
rect 4508 19552 4572 19556
rect 9581 19612 9645 19616
rect 9581 19556 9585 19612
rect 9585 19556 9641 19612
rect 9641 19556 9645 19612
rect 9581 19552 9645 19556
rect 9661 19612 9725 19616
rect 9661 19556 9665 19612
rect 9665 19556 9721 19612
rect 9721 19556 9725 19612
rect 9661 19552 9725 19556
rect 9741 19612 9805 19616
rect 9741 19556 9745 19612
rect 9745 19556 9801 19612
rect 9801 19556 9805 19612
rect 9741 19552 9805 19556
rect 9821 19612 9885 19616
rect 9821 19556 9825 19612
rect 9825 19556 9881 19612
rect 9881 19556 9885 19612
rect 9821 19552 9885 19556
rect 14894 19612 14958 19616
rect 14894 19556 14898 19612
rect 14898 19556 14954 19612
rect 14954 19556 14958 19612
rect 14894 19552 14958 19556
rect 14974 19612 15038 19616
rect 14974 19556 14978 19612
rect 14978 19556 15034 19612
rect 15034 19556 15038 19612
rect 14974 19552 15038 19556
rect 15054 19612 15118 19616
rect 15054 19556 15058 19612
rect 15058 19556 15114 19612
rect 15114 19556 15118 19612
rect 15054 19552 15118 19556
rect 15134 19612 15198 19616
rect 15134 19556 15138 19612
rect 15138 19556 15194 19612
rect 15194 19556 15198 19612
rect 15134 19552 15198 19556
rect 20207 19612 20271 19616
rect 20207 19556 20211 19612
rect 20211 19556 20267 19612
rect 20267 19556 20271 19612
rect 20207 19552 20271 19556
rect 20287 19612 20351 19616
rect 20287 19556 20291 19612
rect 20291 19556 20347 19612
rect 20347 19556 20351 19612
rect 20287 19552 20351 19556
rect 20367 19612 20431 19616
rect 20367 19556 20371 19612
rect 20371 19556 20427 19612
rect 20427 19556 20431 19612
rect 20367 19552 20431 19556
rect 20447 19612 20511 19616
rect 20447 19556 20451 19612
rect 20451 19556 20507 19612
rect 20507 19556 20511 19612
rect 20447 19552 20511 19556
rect 3608 19068 3672 19072
rect 3608 19012 3612 19068
rect 3612 19012 3668 19068
rect 3668 19012 3672 19068
rect 3608 19008 3672 19012
rect 3688 19068 3752 19072
rect 3688 19012 3692 19068
rect 3692 19012 3748 19068
rect 3748 19012 3752 19068
rect 3688 19008 3752 19012
rect 3768 19068 3832 19072
rect 3768 19012 3772 19068
rect 3772 19012 3828 19068
rect 3828 19012 3832 19068
rect 3768 19008 3832 19012
rect 3848 19068 3912 19072
rect 3848 19012 3852 19068
rect 3852 19012 3908 19068
rect 3908 19012 3912 19068
rect 3848 19008 3912 19012
rect 8921 19068 8985 19072
rect 8921 19012 8925 19068
rect 8925 19012 8981 19068
rect 8981 19012 8985 19068
rect 8921 19008 8985 19012
rect 9001 19068 9065 19072
rect 9001 19012 9005 19068
rect 9005 19012 9061 19068
rect 9061 19012 9065 19068
rect 9001 19008 9065 19012
rect 9081 19068 9145 19072
rect 9081 19012 9085 19068
rect 9085 19012 9141 19068
rect 9141 19012 9145 19068
rect 9081 19008 9145 19012
rect 9161 19068 9225 19072
rect 9161 19012 9165 19068
rect 9165 19012 9221 19068
rect 9221 19012 9225 19068
rect 9161 19008 9225 19012
rect 14234 19068 14298 19072
rect 14234 19012 14238 19068
rect 14238 19012 14294 19068
rect 14294 19012 14298 19068
rect 14234 19008 14298 19012
rect 14314 19068 14378 19072
rect 14314 19012 14318 19068
rect 14318 19012 14374 19068
rect 14374 19012 14378 19068
rect 14314 19008 14378 19012
rect 14394 19068 14458 19072
rect 14394 19012 14398 19068
rect 14398 19012 14454 19068
rect 14454 19012 14458 19068
rect 14394 19008 14458 19012
rect 14474 19068 14538 19072
rect 14474 19012 14478 19068
rect 14478 19012 14534 19068
rect 14534 19012 14538 19068
rect 14474 19008 14538 19012
rect 19547 19068 19611 19072
rect 19547 19012 19551 19068
rect 19551 19012 19607 19068
rect 19607 19012 19611 19068
rect 19547 19008 19611 19012
rect 19627 19068 19691 19072
rect 19627 19012 19631 19068
rect 19631 19012 19687 19068
rect 19687 19012 19691 19068
rect 19627 19008 19691 19012
rect 19707 19068 19771 19072
rect 19707 19012 19711 19068
rect 19711 19012 19767 19068
rect 19767 19012 19771 19068
rect 19707 19008 19771 19012
rect 19787 19068 19851 19072
rect 19787 19012 19791 19068
rect 19791 19012 19847 19068
rect 19847 19012 19851 19068
rect 19787 19008 19851 19012
rect 4268 18524 4332 18528
rect 4268 18468 4272 18524
rect 4272 18468 4328 18524
rect 4328 18468 4332 18524
rect 4268 18464 4332 18468
rect 4348 18524 4412 18528
rect 4348 18468 4352 18524
rect 4352 18468 4408 18524
rect 4408 18468 4412 18524
rect 4348 18464 4412 18468
rect 4428 18524 4492 18528
rect 4428 18468 4432 18524
rect 4432 18468 4488 18524
rect 4488 18468 4492 18524
rect 4428 18464 4492 18468
rect 4508 18524 4572 18528
rect 4508 18468 4512 18524
rect 4512 18468 4568 18524
rect 4568 18468 4572 18524
rect 4508 18464 4572 18468
rect 9581 18524 9645 18528
rect 9581 18468 9585 18524
rect 9585 18468 9641 18524
rect 9641 18468 9645 18524
rect 9581 18464 9645 18468
rect 9661 18524 9725 18528
rect 9661 18468 9665 18524
rect 9665 18468 9721 18524
rect 9721 18468 9725 18524
rect 9661 18464 9725 18468
rect 9741 18524 9805 18528
rect 9741 18468 9745 18524
rect 9745 18468 9801 18524
rect 9801 18468 9805 18524
rect 9741 18464 9805 18468
rect 9821 18524 9885 18528
rect 9821 18468 9825 18524
rect 9825 18468 9881 18524
rect 9881 18468 9885 18524
rect 9821 18464 9885 18468
rect 14894 18524 14958 18528
rect 14894 18468 14898 18524
rect 14898 18468 14954 18524
rect 14954 18468 14958 18524
rect 14894 18464 14958 18468
rect 14974 18524 15038 18528
rect 14974 18468 14978 18524
rect 14978 18468 15034 18524
rect 15034 18468 15038 18524
rect 14974 18464 15038 18468
rect 15054 18524 15118 18528
rect 15054 18468 15058 18524
rect 15058 18468 15114 18524
rect 15114 18468 15118 18524
rect 15054 18464 15118 18468
rect 15134 18524 15198 18528
rect 15134 18468 15138 18524
rect 15138 18468 15194 18524
rect 15194 18468 15198 18524
rect 15134 18464 15198 18468
rect 20207 18524 20271 18528
rect 20207 18468 20211 18524
rect 20211 18468 20267 18524
rect 20267 18468 20271 18524
rect 20207 18464 20271 18468
rect 20287 18524 20351 18528
rect 20287 18468 20291 18524
rect 20291 18468 20347 18524
rect 20347 18468 20351 18524
rect 20287 18464 20351 18468
rect 20367 18524 20431 18528
rect 20367 18468 20371 18524
rect 20371 18468 20427 18524
rect 20427 18468 20431 18524
rect 20367 18464 20431 18468
rect 20447 18524 20511 18528
rect 20447 18468 20451 18524
rect 20451 18468 20507 18524
rect 20507 18468 20511 18524
rect 20447 18464 20511 18468
rect 3608 17980 3672 17984
rect 3608 17924 3612 17980
rect 3612 17924 3668 17980
rect 3668 17924 3672 17980
rect 3608 17920 3672 17924
rect 3688 17980 3752 17984
rect 3688 17924 3692 17980
rect 3692 17924 3748 17980
rect 3748 17924 3752 17980
rect 3688 17920 3752 17924
rect 3768 17980 3832 17984
rect 3768 17924 3772 17980
rect 3772 17924 3828 17980
rect 3828 17924 3832 17980
rect 3768 17920 3832 17924
rect 3848 17980 3912 17984
rect 3848 17924 3852 17980
rect 3852 17924 3908 17980
rect 3908 17924 3912 17980
rect 3848 17920 3912 17924
rect 8921 17980 8985 17984
rect 8921 17924 8925 17980
rect 8925 17924 8981 17980
rect 8981 17924 8985 17980
rect 8921 17920 8985 17924
rect 9001 17980 9065 17984
rect 9001 17924 9005 17980
rect 9005 17924 9061 17980
rect 9061 17924 9065 17980
rect 9001 17920 9065 17924
rect 9081 17980 9145 17984
rect 9081 17924 9085 17980
rect 9085 17924 9141 17980
rect 9141 17924 9145 17980
rect 9081 17920 9145 17924
rect 9161 17980 9225 17984
rect 9161 17924 9165 17980
rect 9165 17924 9221 17980
rect 9221 17924 9225 17980
rect 9161 17920 9225 17924
rect 14234 17980 14298 17984
rect 14234 17924 14238 17980
rect 14238 17924 14294 17980
rect 14294 17924 14298 17980
rect 14234 17920 14298 17924
rect 14314 17980 14378 17984
rect 14314 17924 14318 17980
rect 14318 17924 14374 17980
rect 14374 17924 14378 17980
rect 14314 17920 14378 17924
rect 14394 17980 14458 17984
rect 14394 17924 14398 17980
rect 14398 17924 14454 17980
rect 14454 17924 14458 17980
rect 14394 17920 14458 17924
rect 14474 17980 14538 17984
rect 14474 17924 14478 17980
rect 14478 17924 14534 17980
rect 14534 17924 14538 17980
rect 14474 17920 14538 17924
rect 19547 17980 19611 17984
rect 19547 17924 19551 17980
rect 19551 17924 19607 17980
rect 19607 17924 19611 17980
rect 19547 17920 19611 17924
rect 19627 17980 19691 17984
rect 19627 17924 19631 17980
rect 19631 17924 19687 17980
rect 19687 17924 19691 17980
rect 19627 17920 19691 17924
rect 19707 17980 19771 17984
rect 19707 17924 19711 17980
rect 19711 17924 19767 17980
rect 19767 17924 19771 17980
rect 19707 17920 19771 17924
rect 19787 17980 19851 17984
rect 19787 17924 19791 17980
rect 19791 17924 19847 17980
rect 19847 17924 19851 17980
rect 19787 17920 19851 17924
rect 4268 17436 4332 17440
rect 4268 17380 4272 17436
rect 4272 17380 4328 17436
rect 4328 17380 4332 17436
rect 4268 17376 4332 17380
rect 4348 17436 4412 17440
rect 4348 17380 4352 17436
rect 4352 17380 4408 17436
rect 4408 17380 4412 17436
rect 4348 17376 4412 17380
rect 4428 17436 4492 17440
rect 4428 17380 4432 17436
rect 4432 17380 4488 17436
rect 4488 17380 4492 17436
rect 4428 17376 4492 17380
rect 4508 17436 4572 17440
rect 4508 17380 4512 17436
rect 4512 17380 4568 17436
rect 4568 17380 4572 17436
rect 4508 17376 4572 17380
rect 9581 17436 9645 17440
rect 9581 17380 9585 17436
rect 9585 17380 9641 17436
rect 9641 17380 9645 17436
rect 9581 17376 9645 17380
rect 9661 17436 9725 17440
rect 9661 17380 9665 17436
rect 9665 17380 9721 17436
rect 9721 17380 9725 17436
rect 9661 17376 9725 17380
rect 9741 17436 9805 17440
rect 9741 17380 9745 17436
rect 9745 17380 9801 17436
rect 9801 17380 9805 17436
rect 9741 17376 9805 17380
rect 9821 17436 9885 17440
rect 9821 17380 9825 17436
rect 9825 17380 9881 17436
rect 9881 17380 9885 17436
rect 9821 17376 9885 17380
rect 14894 17436 14958 17440
rect 14894 17380 14898 17436
rect 14898 17380 14954 17436
rect 14954 17380 14958 17436
rect 14894 17376 14958 17380
rect 14974 17436 15038 17440
rect 14974 17380 14978 17436
rect 14978 17380 15034 17436
rect 15034 17380 15038 17436
rect 14974 17376 15038 17380
rect 15054 17436 15118 17440
rect 15054 17380 15058 17436
rect 15058 17380 15114 17436
rect 15114 17380 15118 17436
rect 15054 17376 15118 17380
rect 15134 17436 15198 17440
rect 15134 17380 15138 17436
rect 15138 17380 15194 17436
rect 15194 17380 15198 17436
rect 15134 17376 15198 17380
rect 20207 17436 20271 17440
rect 20207 17380 20211 17436
rect 20211 17380 20267 17436
rect 20267 17380 20271 17436
rect 20207 17376 20271 17380
rect 20287 17436 20351 17440
rect 20287 17380 20291 17436
rect 20291 17380 20347 17436
rect 20347 17380 20351 17436
rect 20287 17376 20351 17380
rect 20367 17436 20431 17440
rect 20367 17380 20371 17436
rect 20371 17380 20427 17436
rect 20427 17380 20431 17436
rect 20367 17376 20431 17380
rect 20447 17436 20511 17440
rect 20447 17380 20451 17436
rect 20451 17380 20507 17436
rect 20507 17380 20511 17436
rect 20447 17376 20511 17380
rect 3608 16892 3672 16896
rect 3608 16836 3612 16892
rect 3612 16836 3668 16892
rect 3668 16836 3672 16892
rect 3608 16832 3672 16836
rect 3688 16892 3752 16896
rect 3688 16836 3692 16892
rect 3692 16836 3748 16892
rect 3748 16836 3752 16892
rect 3688 16832 3752 16836
rect 3768 16892 3832 16896
rect 3768 16836 3772 16892
rect 3772 16836 3828 16892
rect 3828 16836 3832 16892
rect 3768 16832 3832 16836
rect 3848 16892 3912 16896
rect 3848 16836 3852 16892
rect 3852 16836 3908 16892
rect 3908 16836 3912 16892
rect 3848 16832 3912 16836
rect 8921 16892 8985 16896
rect 8921 16836 8925 16892
rect 8925 16836 8981 16892
rect 8981 16836 8985 16892
rect 8921 16832 8985 16836
rect 9001 16892 9065 16896
rect 9001 16836 9005 16892
rect 9005 16836 9061 16892
rect 9061 16836 9065 16892
rect 9001 16832 9065 16836
rect 9081 16892 9145 16896
rect 9081 16836 9085 16892
rect 9085 16836 9141 16892
rect 9141 16836 9145 16892
rect 9081 16832 9145 16836
rect 9161 16892 9225 16896
rect 9161 16836 9165 16892
rect 9165 16836 9221 16892
rect 9221 16836 9225 16892
rect 9161 16832 9225 16836
rect 14234 16892 14298 16896
rect 14234 16836 14238 16892
rect 14238 16836 14294 16892
rect 14294 16836 14298 16892
rect 14234 16832 14298 16836
rect 14314 16892 14378 16896
rect 14314 16836 14318 16892
rect 14318 16836 14374 16892
rect 14374 16836 14378 16892
rect 14314 16832 14378 16836
rect 14394 16892 14458 16896
rect 14394 16836 14398 16892
rect 14398 16836 14454 16892
rect 14454 16836 14458 16892
rect 14394 16832 14458 16836
rect 14474 16892 14538 16896
rect 14474 16836 14478 16892
rect 14478 16836 14534 16892
rect 14534 16836 14538 16892
rect 14474 16832 14538 16836
rect 19547 16892 19611 16896
rect 19547 16836 19551 16892
rect 19551 16836 19607 16892
rect 19607 16836 19611 16892
rect 19547 16832 19611 16836
rect 19627 16892 19691 16896
rect 19627 16836 19631 16892
rect 19631 16836 19687 16892
rect 19687 16836 19691 16892
rect 19627 16832 19691 16836
rect 19707 16892 19771 16896
rect 19707 16836 19711 16892
rect 19711 16836 19767 16892
rect 19767 16836 19771 16892
rect 19707 16832 19771 16836
rect 19787 16892 19851 16896
rect 19787 16836 19791 16892
rect 19791 16836 19847 16892
rect 19847 16836 19851 16892
rect 19787 16832 19851 16836
rect 4268 16348 4332 16352
rect 4268 16292 4272 16348
rect 4272 16292 4328 16348
rect 4328 16292 4332 16348
rect 4268 16288 4332 16292
rect 4348 16348 4412 16352
rect 4348 16292 4352 16348
rect 4352 16292 4408 16348
rect 4408 16292 4412 16348
rect 4348 16288 4412 16292
rect 4428 16348 4492 16352
rect 4428 16292 4432 16348
rect 4432 16292 4488 16348
rect 4488 16292 4492 16348
rect 4428 16288 4492 16292
rect 4508 16348 4572 16352
rect 4508 16292 4512 16348
rect 4512 16292 4568 16348
rect 4568 16292 4572 16348
rect 4508 16288 4572 16292
rect 9581 16348 9645 16352
rect 9581 16292 9585 16348
rect 9585 16292 9641 16348
rect 9641 16292 9645 16348
rect 9581 16288 9645 16292
rect 9661 16348 9725 16352
rect 9661 16292 9665 16348
rect 9665 16292 9721 16348
rect 9721 16292 9725 16348
rect 9661 16288 9725 16292
rect 9741 16348 9805 16352
rect 9741 16292 9745 16348
rect 9745 16292 9801 16348
rect 9801 16292 9805 16348
rect 9741 16288 9805 16292
rect 9821 16348 9885 16352
rect 9821 16292 9825 16348
rect 9825 16292 9881 16348
rect 9881 16292 9885 16348
rect 9821 16288 9885 16292
rect 14894 16348 14958 16352
rect 14894 16292 14898 16348
rect 14898 16292 14954 16348
rect 14954 16292 14958 16348
rect 14894 16288 14958 16292
rect 14974 16348 15038 16352
rect 14974 16292 14978 16348
rect 14978 16292 15034 16348
rect 15034 16292 15038 16348
rect 14974 16288 15038 16292
rect 15054 16348 15118 16352
rect 15054 16292 15058 16348
rect 15058 16292 15114 16348
rect 15114 16292 15118 16348
rect 15054 16288 15118 16292
rect 15134 16348 15198 16352
rect 15134 16292 15138 16348
rect 15138 16292 15194 16348
rect 15194 16292 15198 16348
rect 15134 16288 15198 16292
rect 20207 16348 20271 16352
rect 20207 16292 20211 16348
rect 20211 16292 20267 16348
rect 20267 16292 20271 16348
rect 20207 16288 20271 16292
rect 20287 16348 20351 16352
rect 20287 16292 20291 16348
rect 20291 16292 20347 16348
rect 20347 16292 20351 16348
rect 20287 16288 20351 16292
rect 20367 16348 20431 16352
rect 20367 16292 20371 16348
rect 20371 16292 20427 16348
rect 20427 16292 20431 16348
rect 20367 16288 20431 16292
rect 20447 16348 20511 16352
rect 20447 16292 20451 16348
rect 20451 16292 20507 16348
rect 20507 16292 20511 16348
rect 20447 16288 20511 16292
rect 3608 15804 3672 15808
rect 3608 15748 3612 15804
rect 3612 15748 3668 15804
rect 3668 15748 3672 15804
rect 3608 15744 3672 15748
rect 3688 15804 3752 15808
rect 3688 15748 3692 15804
rect 3692 15748 3748 15804
rect 3748 15748 3752 15804
rect 3688 15744 3752 15748
rect 3768 15804 3832 15808
rect 3768 15748 3772 15804
rect 3772 15748 3828 15804
rect 3828 15748 3832 15804
rect 3768 15744 3832 15748
rect 3848 15804 3912 15808
rect 3848 15748 3852 15804
rect 3852 15748 3908 15804
rect 3908 15748 3912 15804
rect 3848 15744 3912 15748
rect 8921 15804 8985 15808
rect 8921 15748 8925 15804
rect 8925 15748 8981 15804
rect 8981 15748 8985 15804
rect 8921 15744 8985 15748
rect 9001 15804 9065 15808
rect 9001 15748 9005 15804
rect 9005 15748 9061 15804
rect 9061 15748 9065 15804
rect 9001 15744 9065 15748
rect 9081 15804 9145 15808
rect 9081 15748 9085 15804
rect 9085 15748 9141 15804
rect 9141 15748 9145 15804
rect 9081 15744 9145 15748
rect 9161 15804 9225 15808
rect 9161 15748 9165 15804
rect 9165 15748 9221 15804
rect 9221 15748 9225 15804
rect 9161 15744 9225 15748
rect 14234 15804 14298 15808
rect 14234 15748 14238 15804
rect 14238 15748 14294 15804
rect 14294 15748 14298 15804
rect 14234 15744 14298 15748
rect 14314 15804 14378 15808
rect 14314 15748 14318 15804
rect 14318 15748 14374 15804
rect 14374 15748 14378 15804
rect 14314 15744 14378 15748
rect 14394 15804 14458 15808
rect 14394 15748 14398 15804
rect 14398 15748 14454 15804
rect 14454 15748 14458 15804
rect 14394 15744 14458 15748
rect 14474 15804 14538 15808
rect 14474 15748 14478 15804
rect 14478 15748 14534 15804
rect 14534 15748 14538 15804
rect 14474 15744 14538 15748
rect 19547 15804 19611 15808
rect 19547 15748 19551 15804
rect 19551 15748 19607 15804
rect 19607 15748 19611 15804
rect 19547 15744 19611 15748
rect 19627 15804 19691 15808
rect 19627 15748 19631 15804
rect 19631 15748 19687 15804
rect 19687 15748 19691 15804
rect 19627 15744 19691 15748
rect 19707 15804 19771 15808
rect 19707 15748 19711 15804
rect 19711 15748 19767 15804
rect 19767 15748 19771 15804
rect 19707 15744 19771 15748
rect 19787 15804 19851 15808
rect 19787 15748 19791 15804
rect 19791 15748 19847 15804
rect 19847 15748 19851 15804
rect 19787 15744 19851 15748
rect 4268 15260 4332 15264
rect 4268 15204 4272 15260
rect 4272 15204 4328 15260
rect 4328 15204 4332 15260
rect 4268 15200 4332 15204
rect 4348 15260 4412 15264
rect 4348 15204 4352 15260
rect 4352 15204 4408 15260
rect 4408 15204 4412 15260
rect 4348 15200 4412 15204
rect 4428 15260 4492 15264
rect 4428 15204 4432 15260
rect 4432 15204 4488 15260
rect 4488 15204 4492 15260
rect 4428 15200 4492 15204
rect 4508 15260 4572 15264
rect 4508 15204 4512 15260
rect 4512 15204 4568 15260
rect 4568 15204 4572 15260
rect 4508 15200 4572 15204
rect 9581 15260 9645 15264
rect 9581 15204 9585 15260
rect 9585 15204 9641 15260
rect 9641 15204 9645 15260
rect 9581 15200 9645 15204
rect 9661 15260 9725 15264
rect 9661 15204 9665 15260
rect 9665 15204 9721 15260
rect 9721 15204 9725 15260
rect 9661 15200 9725 15204
rect 9741 15260 9805 15264
rect 9741 15204 9745 15260
rect 9745 15204 9801 15260
rect 9801 15204 9805 15260
rect 9741 15200 9805 15204
rect 9821 15260 9885 15264
rect 9821 15204 9825 15260
rect 9825 15204 9881 15260
rect 9881 15204 9885 15260
rect 9821 15200 9885 15204
rect 14894 15260 14958 15264
rect 14894 15204 14898 15260
rect 14898 15204 14954 15260
rect 14954 15204 14958 15260
rect 14894 15200 14958 15204
rect 14974 15260 15038 15264
rect 14974 15204 14978 15260
rect 14978 15204 15034 15260
rect 15034 15204 15038 15260
rect 14974 15200 15038 15204
rect 15054 15260 15118 15264
rect 15054 15204 15058 15260
rect 15058 15204 15114 15260
rect 15114 15204 15118 15260
rect 15054 15200 15118 15204
rect 15134 15260 15198 15264
rect 15134 15204 15138 15260
rect 15138 15204 15194 15260
rect 15194 15204 15198 15260
rect 15134 15200 15198 15204
rect 20207 15260 20271 15264
rect 20207 15204 20211 15260
rect 20211 15204 20267 15260
rect 20267 15204 20271 15260
rect 20207 15200 20271 15204
rect 20287 15260 20351 15264
rect 20287 15204 20291 15260
rect 20291 15204 20347 15260
rect 20347 15204 20351 15260
rect 20287 15200 20351 15204
rect 20367 15260 20431 15264
rect 20367 15204 20371 15260
rect 20371 15204 20427 15260
rect 20427 15204 20431 15260
rect 20367 15200 20431 15204
rect 20447 15260 20511 15264
rect 20447 15204 20451 15260
rect 20451 15204 20507 15260
rect 20507 15204 20511 15260
rect 20447 15200 20511 15204
rect 3608 14716 3672 14720
rect 3608 14660 3612 14716
rect 3612 14660 3668 14716
rect 3668 14660 3672 14716
rect 3608 14656 3672 14660
rect 3688 14716 3752 14720
rect 3688 14660 3692 14716
rect 3692 14660 3748 14716
rect 3748 14660 3752 14716
rect 3688 14656 3752 14660
rect 3768 14716 3832 14720
rect 3768 14660 3772 14716
rect 3772 14660 3828 14716
rect 3828 14660 3832 14716
rect 3768 14656 3832 14660
rect 3848 14716 3912 14720
rect 3848 14660 3852 14716
rect 3852 14660 3908 14716
rect 3908 14660 3912 14716
rect 3848 14656 3912 14660
rect 8921 14716 8985 14720
rect 8921 14660 8925 14716
rect 8925 14660 8981 14716
rect 8981 14660 8985 14716
rect 8921 14656 8985 14660
rect 9001 14716 9065 14720
rect 9001 14660 9005 14716
rect 9005 14660 9061 14716
rect 9061 14660 9065 14716
rect 9001 14656 9065 14660
rect 9081 14716 9145 14720
rect 9081 14660 9085 14716
rect 9085 14660 9141 14716
rect 9141 14660 9145 14716
rect 9081 14656 9145 14660
rect 9161 14716 9225 14720
rect 9161 14660 9165 14716
rect 9165 14660 9221 14716
rect 9221 14660 9225 14716
rect 9161 14656 9225 14660
rect 14234 14716 14298 14720
rect 14234 14660 14238 14716
rect 14238 14660 14294 14716
rect 14294 14660 14298 14716
rect 14234 14656 14298 14660
rect 14314 14716 14378 14720
rect 14314 14660 14318 14716
rect 14318 14660 14374 14716
rect 14374 14660 14378 14716
rect 14314 14656 14378 14660
rect 14394 14716 14458 14720
rect 14394 14660 14398 14716
rect 14398 14660 14454 14716
rect 14454 14660 14458 14716
rect 14394 14656 14458 14660
rect 14474 14716 14538 14720
rect 14474 14660 14478 14716
rect 14478 14660 14534 14716
rect 14534 14660 14538 14716
rect 14474 14656 14538 14660
rect 19547 14716 19611 14720
rect 19547 14660 19551 14716
rect 19551 14660 19607 14716
rect 19607 14660 19611 14716
rect 19547 14656 19611 14660
rect 19627 14716 19691 14720
rect 19627 14660 19631 14716
rect 19631 14660 19687 14716
rect 19687 14660 19691 14716
rect 19627 14656 19691 14660
rect 19707 14716 19771 14720
rect 19707 14660 19711 14716
rect 19711 14660 19767 14716
rect 19767 14660 19771 14716
rect 19707 14656 19771 14660
rect 19787 14716 19851 14720
rect 19787 14660 19791 14716
rect 19791 14660 19847 14716
rect 19847 14660 19851 14716
rect 19787 14656 19851 14660
rect 4268 14172 4332 14176
rect 4268 14116 4272 14172
rect 4272 14116 4328 14172
rect 4328 14116 4332 14172
rect 4268 14112 4332 14116
rect 4348 14172 4412 14176
rect 4348 14116 4352 14172
rect 4352 14116 4408 14172
rect 4408 14116 4412 14172
rect 4348 14112 4412 14116
rect 4428 14172 4492 14176
rect 4428 14116 4432 14172
rect 4432 14116 4488 14172
rect 4488 14116 4492 14172
rect 4428 14112 4492 14116
rect 4508 14172 4572 14176
rect 4508 14116 4512 14172
rect 4512 14116 4568 14172
rect 4568 14116 4572 14172
rect 4508 14112 4572 14116
rect 9581 14172 9645 14176
rect 9581 14116 9585 14172
rect 9585 14116 9641 14172
rect 9641 14116 9645 14172
rect 9581 14112 9645 14116
rect 9661 14172 9725 14176
rect 9661 14116 9665 14172
rect 9665 14116 9721 14172
rect 9721 14116 9725 14172
rect 9661 14112 9725 14116
rect 9741 14172 9805 14176
rect 9741 14116 9745 14172
rect 9745 14116 9801 14172
rect 9801 14116 9805 14172
rect 9741 14112 9805 14116
rect 9821 14172 9885 14176
rect 9821 14116 9825 14172
rect 9825 14116 9881 14172
rect 9881 14116 9885 14172
rect 9821 14112 9885 14116
rect 14894 14172 14958 14176
rect 14894 14116 14898 14172
rect 14898 14116 14954 14172
rect 14954 14116 14958 14172
rect 14894 14112 14958 14116
rect 14974 14172 15038 14176
rect 14974 14116 14978 14172
rect 14978 14116 15034 14172
rect 15034 14116 15038 14172
rect 14974 14112 15038 14116
rect 15054 14172 15118 14176
rect 15054 14116 15058 14172
rect 15058 14116 15114 14172
rect 15114 14116 15118 14172
rect 15054 14112 15118 14116
rect 15134 14172 15198 14176
rect 15134 14116 15138 14172
rect 15138 14116 15194 14172
rect 15194 14116 15198 14172
rect 15134 14112 15198 14116
rect 20207 14172 20271 14176
rect 20207 14116 20211 14172
rect 20211 14116 20267 14172
rect 20267 14116 20271 14172
rect 20207 14112 20271 14116
rect 20287 14172 20351 14176
rect 20287 14116 20291 14172
rect 20291 14116 20347 14172
rect 20347 14116 20351 14172
rect 20287 14112 20351 14116
rect 20367 14172 20431 14176
rect 20367 14116 20371 14172
rect 20371 14116 20427 14172
rect 20427 14116 20431 14172
rect 20367 14112 20431 14116
rect 20447 14172 20511 14176
rect 20447 14116 20451 14172
rect 20451 14116 20507 14172
rect 20507 14116 20511 14172
rect 20447 14112 20511 14116
rect 3608 13628 3672 13632
rect 3608 13572 3612 13628
rect 3612 13572 3668 13628
rect 3668 13572 3672 13628
rect 3608 13568 3672 13572
rect 3688 13628 3752 13632
rect 3688 13572 3692 13628
rect 3692 13572 3748 13628
rect 3748 13572 3752 13628
rect 3688 13568 3752 13572
rect 3768 13628 3832 13632
rect 3768 13572 3772 13628
rect 3772 13572 3828 13628
rect 3828 13572 3832 13628
rect 3768 13568 3832 13572
rect 3848 13628 3912 13632
rect 3848 13572 3852 13628
rect 3852 13572 3908 13628
rect 3908 13572 3912 13628
rect 3848 13568 3912 13572
rect 8921 13628 8985 13632
rect 8921 13572 8925 13628
rect 8925 13572 8981 13628
rect 8981 13572 8985 13628
rect 8921 13568 8985 13572
rect 9001 13628 9065 13632
rect 9001 13572 9005 13628
rect 9005 13572 9061 13628
rect 9061 13572 9065 13628
rect 9001 13568 9065 13572
rect 9081 13628 9145 13632
rect 9081 13572 9085 13628
rect 9085 13572 9141 13628
rect 9141 13572 9145 13628
rect 9081 13568 9145 13572
rect 9161 13628 9225 13632
rect 9161 13572 9165 13628
rect 9165 13572 9221 13628
rect 9221 13572 9225 13628
rect 9161 13568 9225 13572
rect 14234 13628 14298 13632
rect 14234 13572 14238 13628
rect 14238 13572 14294 13628
rect 14294 13572 14298 13628
rect 14234 13568 14298 13572
rect 14314 13628 14378 13632
rect 14314 13572 14318 13628
rect 14318 13572 14374 13628
rect 14374 13572 14378 13628
rect 14314 13568 14378 13572
rect 14394 13628 14458 13632
rect 14394 13572 14398 13628
rect 14398 13572 14454 13628
rect 14454 13572 14458 13628
rect 14394 13568 14458 13572
rect 14474 13628 14538 13632
rect 14474 13572 14478 13628
rect 14478 13572 14534 13628
rect 14534 13572 14538 13628
rect 14474 13568 14538 13572
rect 19547 13628 19611 13632
rect 19547 13572 19551 13628
rect 19551 13572 19607 13628
rect 19607 13572 19611 13628
rect 19547 13568 19611 13572
rect 19627 13628 19691 13632
rect 19627 13572 19631 13628
rect 19631 13572 19687 13628
rect 19687 13572 19691 13628
rect 19627 13568 19691 13572
rect 19707 13628 19771 13632
rect 19707 13572 19711 13628
rect 19711 13572 19767 13628
rect 19767 13572 19771 13628
rect 19707 13568 19771 13572
rect 19787 13628 19851 13632
rect 19787 13572 19791 13628
rect 19791 13572 19847 13628
rect 19847 13572 19851 13628
rect 19787 13568 19851 13572
rect 4268 13084 4332 13088
rect 4268 13028 4272 13084
rect 4272 13028 4328 13084
rect 4328 13028 4332 13084
rect 4268 13024 4332 13028
rect 4348 13084 4412 13088
rect 4348 13028 4352 13084
rect 4352 13028 4408 13084
rect 4408 13028 4412 13084
rect 4348 13024 4412 13028
rect 4428 13084 4492 13088
rect 4428 13028 4432 13084
rect 4432 13028 4488 13084
rect 4488 13028 4492 13084
rect 4428 13024 4492 13028
rect 4508 13084 4572 13088
rect 4508 13028 4512 13084
rect 4512 13028 4568 13084
rect 4568 13028 4572 13084
rect 4508 13024 4572 13028
rect 9581 13084 9645 13088
rect 9581 13028 9585 13084
rect 9585 13028 9641 13084
rect 9641 13028 9645 13084
rect 9581 13024 9645 13028
rect 9661 13084 9725 13088
rect 9661 13028 9665 13084
rect 9665 13028 9721 13084
rect 9721 13028 9725 13084
rect 9661 13024 9725 13028
rect 9741 13084 9805 13088
rect 9741 13028 9745 13084
rect 9745 13028 9801 13084
rect 9801 13028 9805 13084
rect 9741 13024 9805 13028
rect 9821 13084 9885 13088
rect 9821 13028 9825 13084
rect 9825 13028 9881 13084
rect 9881 13028 9885 13084
rect 9821 13024 9885 13028
rect 14894 13084 14958 13088
rect 14894 13028 14898 13084
rect 14898 13028 14954 13084
rect 14954 13028 14958 13084
rect 14894 13024 14958 13028
rect 14974 13084 15038 13088
rect 14974 13028 14978 13084
rect 14978 13028 15034 13084
rect 15034 13028 15038 13084
rect 14974 13024 15038 13028
rect 15054 13084 15118 13088
rect 15054 13028 15058 13084
rect 15058 13028 15114 13084
rect 15114 13028 15118 13084
rect 15054 13024 15118 13028
rect 15134 13084 15198 13088
rect 15134 13028 15138 13084
rect 15138 13028 15194 13084
rect 15194 13028 15198 13084
rect 15134 13024 15198 13028
rect 20207 13084 20271 13088
rect 20207 13028 20211 13084
rect 20211 13028 20267 13084
rect 20267 13028 20271 13084
rect 20207 13024 20271 13028
rect 20287 13084 20351 13088
rect 20287 13028 20291 13084
rect 20291 13028 20347 13084
rect 20347 13028 20351 13084
rect 20287 13024 20351 13028
rect 20367 13084 20431 13088
rect 20367 13028 20371 13084
rect 20371 13028 20427 13084
rect 20427 13028 20431 13084
rect 20367 13024 20431 13028
rect 20447 13084 20511 13088
rect 20447 13028 20451 13084
rect 20451 13028 20507 13084
rect 20507 13028 20511 13084
rect 20447 13024 20511 13028
rect 3608 12540 3672 12544
rect 3608 12484 3612 12540
rect 3612 12484 3668 12540
rect 3668 12484 3672 12540
rect 3608 12480 3672 12484
rect 3688 12540 3752 12544
rect 3688 12484 3692 12540
rect 3692 12484 3748 12540
rect 3748 12484 3752 12540
rect 3688 12480 3752 12484
rect 3768 12540 3832 12544
rect 3768 12484 3772 12540
rect 3772 12484 3828 12540
rect 3828 12484 3832 12540
rect 3768 12480 3832 12484
rect 3848 12540 3912 12544
rect 3848 12484 3852 12540
rect 3852 12484 3908 12540
rect 3908 12484 3912 12540
rect 3848 12480 3912 12484
rect 8921 12540 8985 12544
rect 8921 12484 8925 12540
rect 8925 12484 8981 12540
rect 8981 12484 8985 12540
rect 8921 12480 8985 12484
rect 9001 12540 9065 12544
rect 9001 12484 9005 12540
rect 9005 12484 9061 12540
rect 9061 12484 9065 12540
rect 9001 12480 9065 12484
rect 9081 12540 9145 12544
rect 9081 12484 9085 12540
rect 9085 12484 9141 12540
rect 9141 12484 9145 12540
rect 9081 12480 9145 12484
rect 9161 12540 9225 12544
rect 9161 12484 9165 12540
rect 9165 12484 9221 12540
rect 9221 12484 9225 12540
rect 9161 12480 9225 12484
rect 14234 12540 14298 12544
rect 14234 12484 14238 12540
rect 14238 12484 14294 12540
rect 14294 12484 14298 12540
rect 14234 12480 14298 12484
rect 14314 12540 14378 12544
rect 14314 12484 14318 12540
rect 14318 12484 14374 12540
rect 14374 12484 14378 12540
rect 14314 12480 14378 12484
rect 14394 12540 14458 12544
rect 14394 12484 14398 12540
rect 14398 12484 14454 12540
rect 14454 12484 14458 12540
rect 14394 12480 14458 12484
rect 14474 12540 14538 12544
rect 14474 12484 14478 12540
rect 14478 12484 14534 12540
rect 14534 12484 14538 12540
rect 14474 12480 14538 12484
rect 19547 12540 19611 12544
rect 19547 12484 19551 12540
rect 19551 12484 19607 12540
rect 19607 12484 19611 12540
rect 19547 12480 19611 12484
rect 19627 12540 19691 12544
rect 19627 12484 19631 12540
rect 19631 12484 19687 12540
rect 19687 12484 19691 12540
rect 19627 12480 19691 12484
rect 19707 12540 19771 12544
rect 19707 12484 19711 12540
rect 19711 12484 19767 12540
rect 19767 12484 19771 12540
rect 19707 12480 19771 12484
rect 19787 12540 19851 12544
rect 19787 12484 19791 12540
rect 19791 12484 19847 12540
rect 19847 12484 19851 12540
rect 19787 12480 19851 12484
rect 4268 11996 4332 12000
rect 4268 11940 4272 11996
rect 4272 11940 4328 11996
rect 4328 11940 4332 11996
rect 4268 11936 4332 11940
rect 4348 11996 4412 12000
rect 4348 11940 4352 11996
rect 4352 11940 4408 11996
rect 4408 11940 4412 11996
rect 4348 11936 4412 11940
rect 4428 11996 4492 12000
rect 4428 11940 4432 11996
rect 4432 11940 4488 11996
rect 4488 11940 4492 11996
rect 4428 11936 4492 11940
rect 4508 11996 4572 12000
rect 4508 11940 4512 11996
rect 4512 11940 4568 11996
rect 4568 11940 4572 11996
rect 4508 11936 4572 11940
rect 9581 11996 9645 12000
rect 9581 11940 9585 11996
rect 9585 11940 9641 11996
rect 9641 11940 9645 11996
rect 9581 11936 9645 11940
rect 9661 11996 9725 12000
rect 9661 11940 9665 11996
rect 9665 11940 9721 11996
rect 9721 11940 9725 11996
rect 9661 11936 9725 11940
rect 9741 11996 9805 12000
rect 9741 11940 9745 11996
rect 9745 11940 9801 11996
rect 9801 11940 9805 11996
rect 9741 11936 9805 11940
rect 9821 11996 9885 12000
rect 9821 11940 9825 11996
rect 9825 11940 9881 11996
rect 9881 11940 9885 11996
rect 9821 11936 9885 11940
rect 14894 11996 14958 12000
rect 14894 11940 14898 11996
rect 14898 11940 14954 11996
rect 14954 11940 14958 11996
rect 14894 11936 14958 11940
rect 14974 11996 15038 12000
rect 14974 11940 14978 11996
rect 14978 11940 15034 11996
rect 15034 11940 15038 11996
rect 14974 11936 15038 11940
rect 15054 11996 15118 12000
rect 15054 11940 15058 11996
rect 15058 11940 15114 11996
rect 15114 11940 15118 11996
rect 15054 11936 15118 11940
rect 15134 11996 15198 12000
rect 15134 11940 15138 11996
rect 15138 11940 15194 11996
rect 15194 11940 15198 11996
rect 15134 11936 15198 11940
rect 20207 11996 20271 12000
rect 20207 11940 20211 11996
rect 20211 11940 20267 11996
rect 20267 11940 20271 11996
rect 20207 11936 20271 11940
rect 20287 11996 20351 12000
rect 20287 11940 20291 11996
rect 20291 11940 20347 11996
rect 20347 11940 20351 11996
rect 20287 11936 20351 11940
rect 20367 11996 20431 12000
rect 20367 11940 20371 11996
rect 20371 11940 20427 11996
rect 20427 11940 20431 11996
rect 20367 11936 20431 11940
rect 20447 11996 20511 12000
rect 20447 11940 20451 11996
rect 20451 11940 20507 11996
rect 20507 11940 20511 11996
rect 20447 11936 20511 11940
rect 3608 11452 3672 11456
rect 3608 11396 3612 11452
rect 3612 11396 3668 11452
rect 3668 11396 3672 11452
rect 3608 11392 3672 11396
rect 3688 11452 3752 11456
rect 3688 11396 3692 11452
rect 3692 11396 3748 11452
rect 3748 11396 3752 11452
rect 3688 11392 3752 11396
rect 3768 11452 3832 11456
rect 3768 11396 3772 11452
rect 3772 11396 3828 11452
rect 3828 11396 3832 11452
rect 3768 11392 3832 11396
rect 3848 11452 3912 11456
rect 3848 11396 3852 11452
rect 3852 11396 3908 11452
rect 3908 11396 3912 11452
rect 3848 11392 3912 11396
rect 8921 11452 8985 11456
rect 8921 11396 8925 11452
rect 8925 11396 8981 11452
rect 8981 11396 8985 11452
rect 8921 11392 8985 11396
rect 9001 11452 9065 11456
rect 9001 11396 9005 11452
rect 9005 11396 9061 11452
rect 9061 11396 9065 11452
rect 9001 11392 9065 11396
rect 9081 11452 9145 11456
rect 9081 11396 9085 11452
rect 9085 11396 9141 11452
rect 9141 11396 9145 11452
rect 9081 11392 9145 11396
rect 9161 11452 9225 11456
rect 9161 11396 9165 11452
rect 9165 11396 9221 11452
rect 9221 11396 9225 11452
rect 9161 11392 9225 11396
rect 14234 11452 14298 11456
rect 14234 11396 14238 11452
rect 14238 11396 14294 11452
rect 14294 11396 14298 11452
rect 14234 11392 14298 11396
rect 14314 11452 14378 11456
rect 14314 11396 14318 11452
rect 14318 11396 14374 11452
rect 14374 11396 14378 11452
rect 14314 11392 14378 11396
rect 14394 11452 14458 11456
rect 14394 11396 14398 11452
rect 14398 11396 14454 11452
rect 14454 11396 14458 11452
rect 14394 11392 14458 11396
rect 14474 11452 14538 11456
rect 14474 11396 14478 11452
rect 14478 11396 14534 11452
rect 14534 11396 14538 11452
rect 14474 11392 14538 11396
rect 19547 11452 19611 11456
rect 19547 11396 19551 11452
rect 19551 11396 19607 11452
rect 19607 11396 19611 11452
rect 19547 11392 19611 11396
rect 19627 11452 19691 11456
rect 19627 11396 19631 11452
rect 19631 11396 19687 11452
rect 19687 11396 19691 11452
rect 19627 11392 19691 11396
rect 19707 11452 19771 11456
rect 19707 11396 19711 11452
rect 19711 11396 19767 11452
rect 19767 11396 19771 11452
rect 19707 11392 19771 11396
rect 19787 11452 19851 11456
rect 19787 11396 19791 11452
rect 19791 11396 19847 11452
rect 19847 11396 19851 11452
rect 19787 11392 19851 11396
rect 4268 10908 4332 10912
rect 4268 10852 4272 10908
rect 4272 10852 4328 10908
rect 4328 10852 4332 10908
rect 4268 10848 4332 10852
rect 4348 10908 4412 10912
rect 4348 10852 4352 10908
rect 4352 10852 4408 10908
rect 4408 10852 4412 10908
rect 4348 10848 4412 10852
rect 4428 10908 4492 10912
rect 4428 10852 4432 10908
rect 4432 10852 4488 10908
rect 4488 10852 4492 10908
rect 4428 10848 4492 10852
rect 4508 10908 4572 10912
rect 4508 10852 4512 10908
rect 4512 10852 4568 10908
rect 4568 10852 4572 10908
rect 4508 10848 4572 10852
rect 9581 10908 9645 10912
rect 9581 10852 9585 10908
rect 9585 10852 9641 10908
rect 9641 10852 9645 10908
rect 9581 10848 9645 10852
rect 9661 10908 9725 10912
rect 9661 10852 9665 10908
rect 9665 10852 9721 10908
rect 9721 10852 9725 10908
rect 9661 10848 9725 10852
rect 9741 10908 9805 10912
rect 9741 10852 9745 10908
rect 9745 10852 9801 10908
rect 9801 10852 9805 10908
rect 9741 10848 9805 10852
rect 9821 10908 9885 10912
rect 9821 10852 9825 10908
rect 9825 10852 9881 10908
rect 9881 10852 9885 10908
rect 9821 10848 9885 10852
rect 14894 10908 14958 10912
rect 14894 10852 14898 10908
rect 14898 10852 14954 10908
rect 14954 10852 14958 10908
rect 14894 10848 14958 10852
rect 14974 10908 15038 10912
rect 14974 10852 14978 10908
rect 14978 10852 15034 10908
rect 15034 10852 15038 10908
rect 14974 10848 15038 10852
rect 15054 10908 15118 10912
rect 15054 10852 15058 10908
rect 15058 10852 15114 10908
rect 15114 10852 15118 10908
rect 15054 10848 15118 10852
rect 15134 10908 15198 10912
rect 15134 10852 15138 10908
rect 15138 10852 15194 10908
rect 15194 10852 15198 10908
rect 15134 10848 15198 10852
rect 20207 10908 20271 10912
rect 20207 10852 20211 10908
rect 20211 10852 20267 10908
rect 20267 10852 20271 10908
rect 20207 10848 20271 10852
rect 20287 10908 20351 10912
rect 20287 10852 20291 10908
rect 20291 10852 20347 10908
rect 20347 10852 20351 10908
rect 20287 10848 20351 10852
rect 20367 10908 20431 10912
rect 20367 10852 20371 10908
rect 20371 10852 20427 10908
rect 20427 10852 20431 10908
rect 20367 10848 20431 10852
rect 20447 10908 20511 10912
rect 20447 10852 20451 10908
rect 20451 10852 20507 10908
rect 20507 10852 20511 10908
rect 20447 10848 20511 10852
rect 3608 10364 3672 10368
rect 3608 10308 3612 10364
rect 3612 10308 3668 10364
rect 3668 10308 3672 10364
rect 3608 10304 3672 10308
rect 3688 10364 3752 10368
rect 3688 10308 3692 10364
rect 3692 10308 3748 10364
rect 3748 10308 3752 10364
rect 3688 10304 3752 10308
rect 3768 10364 3832 10368
rect 3768 10308 3772 10364
rect 3772 10308 3828 10364
rect 3828 10308 3832 10364
rect 3768 10304 3832 10308
rect 3848 10364 3912 10368
rect 3848 10308 3852 10364
rect 3852 10308 3908 10364
rect 3908 10308 3912 10364
rect 3848 10304 3912 10308
rect 8921 10364 8985 10368
rect 8921 10308 8925 10364
rect 8925 10308 8981 10364
rect 8981 10308 8985 10364
rect 8921 10304 8985 10308
rect 9001 10364 9065 10368
rect 9001 10308 9005 10364
rect 9005 10308 9061 10364
rect 9061 10308 9065 10364
rect 9001 10304 9065 10308
rect 9081 10364 9145 10368
rect 9081 10308 9085 10364
rect 9085 10308 9141 10364
rect 9141 10308 9145 10364
rect 9081 10304 9145 10308
rect 9161 10364 9225 10368
rect 9161 10308 9165 10364
rect 9165 10308 9221 10364
rect 9221 10308 9225 10364
rect 9161 10304 9225 10308
rect 14234 10364 14298 10368
rect 14234 10308 14238 10364
rect 14238 10308 14294 10364
rect 14294 10308 14298 10364
rect 14234 10304 14298 10308
rect 14314 10364 14378 10368
rect 14314 10308 14318 10364
rect 14318 10308 14374 10364
rect 14374 10308 14378 10364
rect 14314 10304 14378 10308
rect 14394 10364 14458 10368
rect 14394 10308 14398 10364
rect 14398 10308 14454 10364
rect 14454 10308 14458 10364
rect 14394 10304 14458 10308
rect 14474 10364 14538 10368
rect 14474 10308 14478 10364
rect 14478 10308 14534 10364
rect 14534 10308 14538 10364
rect 14474 10304 14538 10308
rect 19547 10364 19611 10368
rect 19547 10308 19551 10364
rect 19551 10308 19607 10364
rect 19607 10308 19611 10364
rect 19547 10304 19611 10308
rect 19627 10364 19691 10368
rect 19627 10308 19631 10364
rect 19631 10308 19687 10364
rect 19687 10308 19691 10364
rect 19627 10304 19691 10308
rect 19707 10364 19771 10368
rect 19707 10308 19711 10364
rect 19711 10308 19767 10364
rect 19767 10308 19771 10364
rect 19707 10304 19771 10308
rect 19787 10364 19851 10368
rect 19787 10308 19791 10364
rect 19791 10308 19847 10364
rect 19847 10308 19851 10364
rect 19787 10304 19851 10308
rect 4268 9820 4332 9824
rect 4268 9764 4272 9820
rect 4272 9764 4328 9820
rect 4328 9764 4332 9820
rect 4268 9760 4332 9764
rect 4348 9820 4412 9824
rect 4348 9764 4352 9820
rect 4352 9764 4408 9820
rect 4408 9764 4412 9820
rect 4348 9760 4412 9764
rect 4428 9820 4492 9824
rect 4428 9764 4432 9820
rect 4432 9764 4488 9820
rect 4488 9764 4492 9820
rect 4428 9760 4492 9764
rect 4508 9820 4572 9824
rect 4508 9764 4512 9820
rect 4512 9764 4568 9820
rect 4568 9764 4572 9820
rect 4508 9760 4572 9764
rect 9581 9820 9645 9824
rect 9581 9764 9585 9820
rect 9585 9764 9641 9820
rect 9641 9764 9645 9820
rect 9581 9760 9645 9764
rect 9661 9820 9725 9824
rect 9661 9764 9665 9820
rect 9665 9764 9721 9820
rect 9721 9764 9725 9820
rect 9661 9760 9725 9764
rect 9741 9820 9805 9824
rect 9741 9764 9745 9820
rect 9745 9764 9801 9820
rect 9801 9764 9805 9820
rect 9741 9760 9805 9764
rect 9821 9820 9885 9824
rect 9821 9764 9825 9820
rect 9825 9764 9881 9820
rect 9881 9764 9885 9820
rect 9821 9760 9885 9764
rect 14894 9820 14958 9824
rect 14894 9764 14898 9820
rect 14898 9764 14954 9820
rect 14954 9764 14958 9820
rect 14894 9760 14958 9764
rect 14974 9820 15038 9824
rect 14974 9764 14978 9820
rect 14978 9764 15034 9820
rect 15034 9764 15038 9820
rect 14974 9760 15038 9764
rect 15054 9820 15118 9824
rect 15054 9764 15058 9820
rect 15058 9764 15114 9820
rect 15114 9764 15118 9820
rect 15054 9760 15118 9764
rect 15134 9820 15198 9824
rect 15134 9764 15138 9820
rect 15138 9764 15194 9820
rect 15194 9764 15198 9820
rect 15134 9760 15198 9764
rect 20207 9820 20271 9824
rect 20207 9764 20211 9820
rect 20211 9764 20267 9820
rect 20267 9764 20271 9820
rect 20207 9760 20271 9764
rect 20287 9820 20351 9824
rect 20287 9764 20291 9820
rect 20291 9764 20347 9820
rect 20347 9764 20351 9820
rect 20287 9760 20351 9764
rect 20367 9820 20431 9824
rect 20367 9764 20371 9820
rect 20371 9764 20427 9820
rect 20427 9764 20431 9820
rect 20367 9760 20431 9764
rect 20447 9820 20511 9824
rect 20447 9764 20451 9820
rect 20451 9764 20507 9820
rect 20507 9764 20511 9820
rect 20447 9760 20511 9764
rect 3608 9276 3672 9280
rect 3608 9220 3612 9276
rect 3612 9220 3668 9276
rect 3668 9220 3672 9276
rect 3608 9216 3672 9220
rect 3688 9276 3752 9280
rect 3688 9220 3692 9276
rect 3692 9220 3748 9276
rect 3748 9220 3752 9276
rect 3688 9216 3752 9220
rect 3768 9276 3832 9280
rect 3768 9220 3772 9276
rect 3772 9220 3828 9276
rect 3828 9220 3832 9276
rect 3768 9216 3832 9220
rect 3848 9276 3912 9280
rect 3848 9220 3852 9276
rect 3852 9220 3908 9276
rect 3908 9220 3912 9276
rect 3848 9216 3912 9220
rect 8921 9276 8985 9280
rect 8921 9220 8925 9276
rect 8925 9220 8981 9276
rect 8981 9220 8985 9276
rect 8921 9216 8985 9220
rect 9001 9276 9065 9280
rect 9001 9220 9005 9276
rect 9005 9220 9061 9276
rect 9061 9220 9065 9276
rect 9001 9216 9065 9220
rect 9081 9276 9145 9280
rect 9081 9220 9085 9276
rect 9085 9220 9141 9276
rect 9141 9220 9145 9276
rect 9081 9216 9145 9220
rect 9161 9276 9225 9280
rect 9161 9220 9165 9276
rect 9165 9220 9221 9276
rect 9221 9220 9225 9276
rect 9161 9216 9225 9220
rect 14234 9276 14298 9280
rect 14234 9220 14238 9276
rect 14238 9220 14294 9276
rect 14294 9220 14298 9276
rect 14234 9216 14298 9220
rect 14314 9276 14378 9280
rect 14314 9220 14318 9276
rect 14318 9220 14374 9276
rect 14374 9220 14378 9276
rect 14314 9216 14378 9220
rect 14394 9276 14458 9280
rect 14394 9220 14398 9276
rect 14398 9220 14454 9276
rect 14454 9220 14458 9276
rect 14394 9216 14458 9220
rect 14474 9276 14538 9280
rect 14474 9220 14478 9276
rect 14478 9220 14534 9276
rect 14534 9220 14538 9276
rect 14474 9216 14538 9220
rect 19547 9276 19611 9280
rect 19547 9220 19551 9276
rect 19551 9220 19607 9276
rect 19607 9220 19611 9276
rect 19547 9216 19611 9220
rect 19627 9276 19691 9280
rect 19627 9220 19631 9276
rect 19631 9220 19687 9276
rect 19687 9220 19691 9276
rect 19627 9216 19691 9220
rect 19707 9276 19771 9280
rect 19707 9220 19711 9276
rect 19711 9220 19767 9276
rect 19767 9220 19771 9276
rect 19707 9216 19771 9220
rect 19787 9276 19851 9280
rect 19787 9220 19791 9276
rect 19791 9220 19847 9276
rect 19847 9220 19851 9276
rect 19787 9216 19851 9220
rect 4268 8732 4332 8736
rect 4268 8676 4272 8732
rect 4272 8676 4328 8732
rect 4328 8676 4332 8732
rect 4268 8672 4332 8676
rect 4348 8732 4412 8736
rect 4348 8676 4352 8732
rect 4352 8676 4408 8732
rect 4408 8676 4412 8732
rect 4348 8672 4412 8676
rect 4428 8732 4492 8736
rect 4428 8676 4432 8732
rect 4432 8676 4488 8732
rect 4488 8676 4492 8732
rect 4428 8672 4492 8676
rect 4508 8732 4572 8736
rect 4508 8676 4512 8732
rect 4512 8676 4568 8732
rect 4568 8676 4572 8732
rect 4508 8672 4572 8676
rect 9581 8732 9645 8736
rect 9581 8676 9585 8732
rect 9585 8676 9641 8732
rect 9641 8676 9645 8732
rect 9581 8672 9645 8676
rect 9661 8732 9725 8736
rect 9661 8676 9665 8732
rect 9665 8676 9721 8732
rect 9721 8676 9725 8732
rect 9661 8672 9725 8676
rect 9741 8732 9805 8736
rect 9741 8676 9745 8732
rect 9745 8676 9801 8732
rect 9801 8676 9805 8732
rect 9741 8672 9805 8676
rect 9821 8732 9885 8736
rect 9821 8676 9825 8732
rect 9825 8676 9881 8732
rect 9881 8676 9885 8732
rect 9821 8672 9885 8676
rect 14894 8732 14958 8736
rect 14894 8676 14898 8732
rect 14898 8676 14954 8732
rect 14954 8676 14958 8732
rect 14894 8672 14958 8676
rect 14974 8732 15038 8736
rect 14974 8676 14978 8732
rect 14978 8676 15034 8732
rect 15034 8676 15038 8732
rect 14974 8672 15038 8676
rect 15054 8732 15118 8736
rect 15054 8676 15058 8732
rect 15058 8676 15114 8732
rect 15114 8676 15118 8732
rect 15054 8672 15118 8676
rect 15134 8732 15198 8736
rect 15134 8676 15138 8732
rect 15138 8676 15194 8732
rect 15194 8676 15198 8732
rect 15134 8672 15198 8676
rect 20207 8732 20271 8736
rect 20207 8676 20211 8732
rect 20211 8676 20267 8732
rect 20267 8676 20271 8732
rect 20207 8672 20271 8676
rect 20287 8732 20351 8736
rect 20287 8676 20291 8732
rect 20291 8676 20347 8732
rect 20347 8676 20351 8732
rect 20287 8672 20351 8676
rect 20367 8732 20431 8736
rect 20367 8676 20371 8732
rect 20371 8676 20427 8732
rect 20427 8676 20431 8732
rect 20367 8672 20431 8676
rect 20447 8732 20511 8736
rect 20447 8676 20451 8732
rect 20451 8676 20507 8732
rect 20507 8676 20511 8732
rect 20447 8672 20511 8676
rect 3608 8188 3672 8192
rect 3608 8132 3612 8188
rect 3612 8132 3668 8188
rect 3668 8132 3672 8188
rect 3608 8128 3672 8132
rect 3688 8188 3752 8192
rect 3688 8132 3692 8188
rect 3692 8132 3748 8188
rect 3748 8132 3752 8188
rect 3688 8128 3752 8132
rect 3768 8188 3832 8192
rect 3768 8132 3772 8188
rect 3772 8132 3828 8188
rect 3828 8132 3832 8188
rect 3768 8128 3832 8132
rect 3848 8188 3912 8192
rect 3848 8132 3852 8188
rect 3852 8132 3908 8188
rect 3908 8132 3912 8188
rect 3848 8128 3912 8132
rect 8921 8188 8985 8192
rect 8921 8132 8925 8188
rect 8925 8132 8981 8188
rect 8981 8132 8985 8188
rect 8921 8128 8985 8132
rect 9001 8188 9065 8192
rect 9001 8132 9005 8188
rect 9005 8132 9061 8188
rect 9061 8132 9065 8188
rect 9001 8128 9065 8132
rect 9081 8188 9145 8192
rect 9081 8132 9085 8188
rect 9085 8132 9141 8188
rect 9141 8132 9145 8188
rect 9081 8128 9145 8132
rect 9161 8188 9225 8192
rect 9161 8132 9165 8188
rect 9165 8132 9221 8188
rect 9221 8132 9225 8188
rect 9161 8128 9225 8132
rect 14234 8188 14298 8192
rect 14234 8132 14238 8188
rect 14238 8132 14294 8188
rect 14294 8132 14298 8188
rect 14234 8128 14298 8132
rect 14314 8188 14378 8192
rect 14314 8132 14318 8188
rect 14318 8132 14374 8188
rect 14374 8132 14378 8188
rect 14314 8128 14378 8132
rect 14394 8188 14458 8192
rect 14394 8132 14398 8188
rect 14398 8132 14454 8188
rect 14454 8132 14458 8188
rect 14394 8128 14458 8132
rect 14474 8188 14538 8192
rect 14474 8132 14478 8188
rect 14478 8132 14534 8188
rect 14534 8132 14538 8188
rect 14474 8128 14538 8132
rect 19547 8188 19611 8192
rect 19547 8132 19551 8188
rect 19551 8132 19607 8188
rect 19607 8132 19611 8188
rect 19547 8128 19611 8132
rect 19627 8188 19691 8192
rect 19627 8132 19631 8188
rect 19631 8132 19687 8188
rect 19687 8132 19691 8188
rect 19627 8128 19691 8132
rect 19707 8188 19771 8192
rect 19707 8132 19711 8188
rect 19711 8132 19767 8188
rect 19767 8132 19771 8188
rect 19707 8128 19771 8132
rect 19787 8188 19851 8192
rect 19787 8132 19791 8188
rect 19791 8132 19847 8188
rect 19847 8132 19851 8188
rect 19787 8128 19851 8132
rect 4268 7644 4332 7648
rect 4268 7588 4272 7644
rect 4272 7588 4328 7644
rect 4328 7588 4332 7644
rect 4268 7584 4332 7588
rect 4348 7644 4412 7648
rect 4348 7588 4352 7644
rect 4352 7588 4408 7644
rect 4408 7588 4412 7644
rect 4348 7584 4412 7588
rect 4428 7644 4492 7648
rect 4428 7588 4432 7644
rect 4432 7588 4488 7644
rect 4488 7588 4492 7644
rect 4428 7584 4492 7588
rect 4508 7644 4572 7648
rect 4508 7588 4512 7644
rect 4512 7588 4568 7644
rect 4568 7588 4572 7644
rect 4508 7584 4572 7588
rect 9581 7644 9645 7648
rect 9581 7588 9585 7644
rect 9585 7588 9641 7644
rect 9641 7588 9645 7644
rect 9581 7584 9645 7588
rect 9661 7644 9725 7648
rect 9661 7588 9665 7644
rect 9665 7588 9721 7644
rect 9721 7588 9725 7644
rect 9661 7584 9725 7588
rect 9741 7644 9805 7648
rect 9741 7588 9745 7644
rect 9745 7588 9801 7644
rect 9801 7588 9805 7644
rect 9741 7584 9805 7588
rect 9821 7644 9885 7648
rect 9821 7588 9825 7644
rect 9825 7588 9881 7644
rect 9881 7588 9885 7644
rect 9821 7584 9885 7588
rect 14894 7644 14958 7648
rect 14894 7588 14898 7644
rect 14898 7588 14954 7644
rect 14954 7588 14958 7644
rect 14894 7584 14958 7588
rect 14974 7644 15038 7648
rect 14974 7588 14978 7644
rect 14978 7588 15034 7644
rect 15034 7588 15038 7644
rect 14974 7584 15038 7588
rect 15054 7644 15118 7648
rect 15054 7588 15058 7644
rect 15058 7588 15114 7644
rect 15114 7588 15118 7644
rect 15054 7584 15118 7588
rect 15134 7644 15198 7648
rect 15134 7588 15138 7644
rect 15138 7588 15194 7644
rect 15194 7588 15198 7644
rect 15134 7584 15198 7588
rect 20207 7644 20271 7648
rect 20207 7588 20211 7644
rect 20211 7588 20267 7644
rect 20267 7588 20271 7644
rect 20207 7584 20271 7588
rect 20287 7644 20351 7648
rect 20287 7588 20291 7644
rect 20291 7588 20347 7644
rect 20347 7588 20351 7644
rect 20287 7584 20351 7588
rect 20367 7644 20431 7648
rect 20367 7588 20371 7644
rect 20371 7588 20427 7644
rect 20427 7588 20431 7644
rect 20367 7584 20431 7588
rect 20447 7644 20511 7648
rect 20447 7588 20451 7644
rect 20451 7588 20507 7644
rect 20507 7588 20511 7644
rect 20447 7584 20511 7588
rect 3608 7100 3672 7104
rect 3608 7044 3612 7100
rect 3612 7044 3668 7100
rect 3668 7044 3672 7100
rect 3608 7040 3672 7044
rect 3688 7100 3752 7104
rect 3688 7044 3692 7100
rect 3692 7044 3748 7100
rect 3748 7044 3752 7100
rect 3688 7040 3752 7044
rect 3768 7100 3832 7104
rect 3768 7044 3772 7100
rect 3772 7044 3828 7100
rect 3828 7044 3832 7100
rect 3768 7040 3832 7044
rect 3848 7100 3912 7104
rect 3848 7044 3852 7100
rect 3852 7044 3908 7100
rect 3908 7044 3912 7100
rect 3848 7040 3912 7044
rect 8921 7100 8985 7104
rect 8921 7044 8925 7100
rect 8925 7044 8981 7100
rect 8981 7044 8985 7100
rect 8921 7040 8985 7044
rect 9001 7100 9065 7104
rect 9001 7044 9005 7100
rect 9005 7044 9061 7100
rect 9061 7044 9065 7100
rect 9001 7040 9065 7044
rect 9081 7100 9145 7104
rect 9081 7044 9085 7100
rect 9085 7044 9141 7100
rect 9141 7044 9145 7100
rect 9081 7040 9145 7044
rect 9161 7100 9225 7104
rect 9161 7044 9165 7100
rect 9165 7044 9221 7100
rect 9221 7044 9225 7100
rect 9161 7040 9225 7044
rect 14234 7100 14298 7104
rect 14234 7044 14238 7100
rect 14238 7044 14294 7100
rect 14294 7044 14298 7100
rect 14234 7040 14298 7044
rect 14314 7100 14378 7104
rect 14314 7044 14318 7100
rect 14318 7044 14374 7100
rect 14374 7044 14378 7100
rect 14314 7040 14378 7044
rect 14394 7100 14458 7104
rect 14394 7044 14398 7100
rect 14398 7044 14454 7100
rect 14454 7044 14458 7100
rect 14394 7040 14458 7044
rect 14474 7100 14538 7104
rect 14474 7044 14478 7100
rect 14478 7044 14534 7100
rect 14534 7044 14538 7100
rect 14474 7040 14538 7044
rect 19547 7100 19611 7104
rect 19547 7044 19551 7100
rect 19551 7044 19607 7100
rect 19607 7044 19611 7100
rect 19547 7040 19611 7044
rect 19627 7100 19691 7104
rect 19627 7044 19631 7100
rect 19631 7044 19687 7100
rect 19687 7044 19691 7100
rect 19627 7040 19691 7044
rect 19707 7100 19771 7104
rect 19707 7044 19711 7100
rect 19711 7044 19767 7100
rect 19767 7044 19771 7100
rect 19707 7040 19771 7044
rect 19787 7100 19851 7104
rect 19787 7044 19791 7100
rect 19791 7044 19847 7100
rect 19847 7044 19851 7100
rect 19787 7040 19851 7044
rect 4268 6556 4332 6560
rect 4268 6500 4272 6556
rect 4272 6500 4328 6556
rect 4328 6500 4332 6556
rect 4268 6496 4332 6500
rect 4348 6556 4412 6560
rect 4348 6500 4352 6556
rect 4352 6500 4408 6556
rect 4408 6500 4412 6556
rect 4348 6496 4412 6500
rect 4428 6556 4492 6560
rect 4428 6500 4432 6556
rect 4432 6500 4488 6556
rect 4488 6500 4492 6556
rect 4428 6496 4492 6500
rect 4508 6556 4572 6560
rect 4508 6500 4512 6556
rect 4512 6500 4568 6556
rect 4568 6500 4572 6556
rect 4508 6496 4572 6500
rect 9581 6556 9645 6560
rect 9581 6500 9585 6556
rect 9585 6500 9641 6556
rect 9641 6500 9645 6556
rect 9581 6496 9645 6500
rect 9661 6556 9725 6560
rect 9661 6500 9665 6556
rect 9665 6500 9721 6556
rect 9721 6500 9725 6556
rect 9661 6496 9725 6500
rect 9741 6556 9805 6560
rect 9741 6500 9745 6556
rect 9745 6500 9801 6556
rect 9801 6500 9805 6556
rect 9741 6496 9805 6500
rect 9821 6556 9885 6560
rect 9821 6500 9825 6556
rect 9825 6500 9881 6556
rect 9881 6500 9885 6556
rect 9821 6496 9885 6500
rect 14894 6556 14958 6560
rect 14894 6500 14898 6556
rect 14898 6500 14954 6556
rect 14954 6500 14958 6556
rect 14894 6496 14958 6500
rect 14974 6556 15038 6560
rect 14974 6500 14978 6556
rect 14978 6500 15034 6556
rect 15034 6500 15038 6556
rect 14974 6496 15038 6500
rect 15054 6556 15118 6560
rect 15054 6500 15058 6556
rect 15058 6500 15114 6556
rect 15114 6500 15118 6556
rect 15054 6496 15118 6500
rect 15134 6556 15198 6560
rect 15134 6500 15138 6556
rect 15138 6500 15194 6556
rect 15194 6500 15198 6556
rect 15134 6496 15198 6500
rect 20207 6556 20271 6560
rect 20207 6500 20211 6556
rect 20211 6500 20267 6556
rect 20267 6500 20271 6556
rect 20207 6496 20271 6500
rect 20287 6556 20351 6560
rect 20287 6500 20291 6556
rect 20291 6500 20347 6556
rect 20347 6500 20351 6556
rect 20287 6496 20351 6500
rect 20367 6556 20431 6560
rect 20367 6500 20371 6556
rect 20371 6500 20427 6556
rect 20427 6500 20431 6556
rect 20367 6496 20431 6500
rect 20447 6556 20511 6560
rect 20447 6500 20451 6556
rect 20451 6500 20507 6556
rect 20507 6500 20511 6556
rect 20447 6496 20511 6500
rect 3608 6012 3672 6016
rect 3608 5956 3612 6012
rect 3612 5956 3668 6012
rect 3668 5956 3672 6012
rect 3608 5952 3672 5956
rect 3688 6012 3752 6016
rect 3688 5956 3692 6012
rect 3692 5956 3748 6012
rect 3748 5956 3752 6012
rect 3688 5952 3752 5956
rect 3768 6012 3832 6016
rect 3768 5956 3772 6012
rect 3772 5956 3828 6012
rect 3828 5956 3832 6012
rect 3768 5952 3832 5956
rect 3848 6012 3912 6016
rect 3848 5956 3852 6012
rect 3852 5956 3908 6012
rect 3908 5956 3912 6012
rect 3848 5952 3912 5956
rect 8921 6012 8985 6016
rect 8921 5956 8925 6012
rect 8925 5956 8981 6012
rect 8981 5956 8985 6012
rect 8921 5952 8985 5956
rect 9001 6012 9065 6016
rect 9001 5956 9005 6012
rect 9005 5956 9061 6012
rect 9061 5956 9065 6012
rect 9001 5952 9065 5956
rect 9081 6012 9145 6016
rect 9081 5956 9085 6012
rect 9085 5956 9141 6012
rect 9141 5956 9145 6012
rect 9081 5952 9145 5956
rect 9161 6012 9225 6016
rect 9161 5956 9165 6012
rect 9165 5956 9221 6012
rect 9221 5956 9225 6012
rect 9161 5952 9225 5956
rect 14234 6012 14298 6016
rect 14234 5956 14238 6012
rect 14238 5956 14294 6012
rect 14294 5956 14298 6012
rect 14234 5952 14298 5956
rect 14314 6012 14378 6016
rect 14314 5956 14318 6012
rect 14318 5956 14374 6012
rect 14374 5956 14378 6012
rect 14314 5952 14378 5956
rect 14394 6012 14458 6016
rect 14394 5956 14398 6012
rect 14398 5956 14454 6012
rect 14454 5956 14458 6012
rect 14394 5952 14458 5956
rect 14474 6012 14538 6016
rect 14474 5956 14478 6012
rect 14478 5956 14534 6012
rect 14534 5956 14538 6012
rect 14474 5952 14538 5956
rect 19547 6012 19611 6016
rect 19547 5956 19551 6012
rect 19551 5956 19607 6012
rect 19607 5956 19611 6012
rect 19547 5952 19611 5956
rect 19627 6012 19691 6016
rect 19627 5956 19631 6012
rect 19631 5956 19687 6012
rect 19687 5956 19691 6012
rect 19627 5952 19691 5956
rect 19707 6012 19771 6016
rect 19707 5956 19711 6012
rect 19711 5956 19767 6012
rect 19767 5956 19771 6012
rect 19707 5952 19771 5956
rect 19787 6012 19851 6016
rect 19787 5956 19791 6012
rect 19791 5956 19847 6012
rect 19847 5956 19851 6012
rect 19787 5952 19851 5956
rect 4268 5468 4332 5472
rect 4268 5412 4272 5468
rect 4272 5412 4328 5468
rect 4328 5412 4332 5468
rect 4268 5408 4332 5412
rect 4348 5468 4412 5472
rect 4348 5412 4352 5468
rect 4352 5412 4408 5468
rect 4408 5412 4412 5468
rect 4348 5408 4412 5412
rect 4428 5468 4492 5472
rect 4428 5412 4432 5468
rect 4432 5412 4488 5468
rect 4488 5412 4492 5468
rect 4428 5408 4492 5412
rect 4508 5468 4572 5472
rect 4508 5412 4512 5468
rect 4512 5412 4568 5468
rect 4568 5412 4572 5468
rect 4508 5408 4572 5412
rect 9581 5468 9645 5472
rect 9581 5412 9585 5468
rect 9585 5412 9641 5468
rect 9641 5412 9645 5468
rect 9581 5408 9645 5412
rect 9661 5468 9725 5472
rect 9661 5412 9665 5468
rect 9665 5412 9721 5468
rect 9721 5412 9725 5468
rect 9661 5408 9725 5412
rect 9741 5468 9805 5472
rect 9741 5412 9745 5468
rect 9745 5412 9801 5468
rect 9801 5412 9805 5468
rect 9741 5408 9805 5412
rect 9821 5468 9885 5472
rect 9821 5412 9825 5468
rect 9825 5412 9881 5468
rect 9881 5412 9885 5468
rect 9821 5408 9885 5412
rect 14894 5468 14958 5472
rect 14894 5412 14898 5468
rect 14898 5412 14954 5468
rect 14954 5412 14958 5468
rect 14894 5408 14958 5412
rect 14974 5468 15038 5472
rect 14974 5412 14978 5468
rect 14978 5412 15034 5468
rect 15034 5412 15038 5468
rect 14974 5408 15038 5412
rect 15054 5468 15118 5472
rect 15054 5412 15058 5468
rect 15058 5412 15114 5468
rect 15114 5412 15118 5468
rect 15054 5408 15118 5412
rect 15134 5468 15198 5472
rect 15134 5412 15138 5468
rect 15138 5412 15194 5468
rect 15194 5412 15198 5468
rect 15134 5408 15198 5412
rect 20207 5468 20271 5472
rect 20207 5412 20211 5468
rect 20211 5412 20267 5468
rect 20267 5412 20271 5468
rect 20207 5408 20271 5412
rect 20287 5468 20351 5472
rect 20287 5412 20291 5468
rect 20291 5412 20347 5468
rect 20347 5412 20351 5468
rect 20287 5408 20351 5412
rect 20367 5468 20431 5472
rect 20367 5412 20371 5468
rect 20371 5412 20427 5468
rect 20427 5412 20431 5468
rect 20367 5408 20431 5412
rect 20447 5468 20511 5472
rect 20447 5412 20451 5468
rect 20451 5412 20507 5468
rect 20507 5412 20511 5468
rect 20447 5408 20511 5412
rect 3608 4924 3672 4928
rect 3608 4868 3612 4924
rect 3612 4868 3668 4924
rect 3668 4868 3672 4924
rect 3608 4864 3672 4868
rect 3688 4924 3752 4928
rect 3688 4868 3692 4924
rect 3692 4868 3748 4924
rect 3748 4868 3752 4924
rect 3688 4864 3752 4868
rect 3768 4924 3832 4928
rect 3768 4868 3772 4924
rect 3772 4868 3828 4924
rect 3828 4868 3832 4924
rect 3768 4864 3832 4868
rect 3848 4924 3912 4928
rect 3848 4868 3852 4924
rect 3852 4868 3908 4924
rect 3908 4868 3912 4924
rect 3848 4864 3912 4868
rect 8921 4924 8985 4928
rect 8921 4868 8925 4924
rect 8925 4868 8981 4924
rect 8981 4868 8985 4924
rect 8921 4864 8985 4868
rect 9001 4924 9065 4928
rect 9001 4868 9005 4924
rect 9005 4868 9061 4924
rect 9061 4868 9065 4924
rect 9001 4864 9065 4868
rect 9081 4924 9145 4928
rect 9081 4868 9085 4924
rect 9085 4868 9141 4924
rect 9141 4868 9145 4924
rect 9081 4864 9145 4868
rect 9161 4924 9225 4928
rect 9161 4868 9165 4924
rect 9165 4868 9221 4924
rect 9221 4868 9225 4924
rect 9161 4864 9225 4868
rect 14234 4924 14298 4928
rect 14234 4868 14238 4924
rect 14238 4868 14294 4924
rect 14294 4868 14298 4924
rect 14234 4864 14298 4868
rect 14314 4924 14378 4928
rect 14314 4868 14318 4924
rect 14318 4868 14374 4924
rect 14374 4868 14378 4924
rect 14314 4864 14378 4868
rect 14394 4924 14458 4928
rect 14394 4868 14398 4924
rect 14398 4868 14454 4924
rect 14454 4868 14458 4924
rect 14394 4864 14458 4868
rect 14474 4924 14538 4928
rect 14474 4868 14478 4924
rect 14478 4868 14534 4924
rect 14534 4868 14538 4924
rect 14474 4864 14538 4868
rect 19547 4924 19611 4928
rect 19547 4868 19551 4924
rect 19551 4868 19607 4924
rect 19607 4868 19611 4924
rect 19547 4864 19611 4868
rect 19627 4924 19691 4928
rect 19627 4868 19631 4924
rect 19631 4868 19687 4924
rect 19687 4868 19691 4924
rect 19627 4864 19691 4868
rect 19707 4924 19771 4928
rect 19707 4868 19711 4924
rect 19711 4868 19767 4924
rect 19767 4868 19771 4924
rect 19707 4864 19771 4868
rect 19787 4924 19851 4928
rect 19787 4868 19791 4924
rect 19791 4868 19847 4924
rect 19847 4868 19851 4924
rect 19787 4864 19851 4868
rect 4268 4380 4332 4384
rect 4268 4324 4272 4380
rect 4272 4324 4328 4380
rect 4328 4324 4332 4380
rect 4268 4320 4332 4324
rect 4348 4380 4412 4384
rect 4348 4324 4352 4380
rect 4352 4324 4408 4380
rect 4408 4324 4412 4380
rect 4348 4320 4412 4324
rect 4428 4380 4492 4384
rect 4428 4324 4432 4380
rect 4432 4324 4488 4380
rect 4488 4324 4492 4380
rect 4428 4320 4492 4324
rect 4508 4380 4572 4384
rect 4508 4324 4512 4380
rect 4512 4324 4568 4380
rect 4568 4324 4572 4380
rect 4508 4320 4572 4324
rect 9581 4380 9645 4384
rect 9581 4324 9585 4380
rect 9585 4324 9641 4380
rect 9641 4324 9645 4380
rect 9581 4320 9645 4324
rect 9661 4380 9725 4384
rect 9661 4324 9665 4380
rect 9665 4324 9721 4380
rect 9721 4324 9725 4380
rect 9661 4320 9725 4324
rect 9741 4380 9805 4384
rect 9741 4324 9745 4380
rect 9745 4324 9801 4380
rect 9801 4324 9805 4380
rect 9741 4320 9805 4324
rect 9821 4380 9885 4384
rect 9821 4324 9825 4380
rect 9825 4324 9881 4380
rect 9881 4324 9885 4380
rect 9821 4320 9885 4324
rect 14894 4380 14958 4384
rect 14894 4324 14898 4380
rect 14898 4324 14954 4380
rect 14954 4324 14958 4380
rect 14894 4320 14958 4324
rect 14974 4380 15038 4384
rect 14974 4324 14978 4380
rect 14978 4324 15034 4380
rect 15034 4324 15038 4380
rect 14974 4320 15038 4324
rect 15054 4380 15118 4384
rect 15054 4324 15058 4380
rect 15058 4324 15114 4380
rect 15114 4324 15118 4380
rect 15054 4320 15118 4324
rect 15134 4380 15198 4384
rect 15134 4324 15138 4380
rect 15138 4324 15194 4380
rect 15194 4324 15198 4380
rect 15134 4320 15198 4324
rect 20207 4380 20271 4384
rect 20207 4324 20211 4380
rect 20211 4324 20267 4380
rect 20267 4324 20271 4380
rect 20207 4320 20271 4324
rect 20287 4380 20351 4384
rect 20287 4324 20291 4380
rect 20291 4324 20347 4380
rect 20347 4324 20351 4380
rect 20287 4320 20351 4324
rect 20367 4380 20431 4384
rect 20367 4324 20371 4380
rect 20371 4324 20427 4380
rect 20427 4324 20431 4380
rect 20367 4320 20431 4324
rect 20447 4380 20511 4384
rect 20447 4324 20451 4380
rect 20451 4324 20507 4380
rect 20507 4324 20511 4380
rect 20447 4320 20511 4324
rect 3608 3836 3672 3840
rect 3608 3780 3612 3836
rect 3612 3780 3668 3836
rect 3668 3780 3672 3836
rect 3608 3776 3672 3780
rect 3688 3836 3752 3840
rect 3688 3780 3692 3836
rect 3692 3780 3748 3836
rect 3748 3780 3752 3836
rect 3688 3776 3752 3780
rect 3768 3836 3832 3840
rect 3768 3780 3772 3836
rect 3772 3780 3828 3836
rect 3828 3780 3832 3836
rect 3768 3776 3832 3780
rect 3848 3836 3912 3840
rect 3848 3780 3852 3836
rect 3852 3780 3908 3836
rect 3908 3780 3912 3836
rect 3848 3776 3912 3780
rect 8921 3836 8985 3840
rect 8921 3780 8925 3836
rect 8925 3780 8981 3836
rect 8981 3780 8985 3836
rect 8921 3776 8985 3780
rect 9001 3836 9065 3840
rect 9001 3780 9005 3836
rect 9005 3780 9061 3836
rect 9061 3780 9065 3836
rect 9001 3776 9065 3780
rect 9081 3836 9145 3840
rect 9081 3780 9085 3836
rect 9085 3780 9141 3836
rect 9141 3780 9145 3836
rect 9081 3776 9145 3780
rect 9161 3836 9225 3840
rect 9161 3780 9165 3836
rect 9165 3780 9221 3836
rect 9221 3780 9225 3836
rect 9161 3776 9225 3780
rect 14234 3836 14298 3840
rect 14234 3780 14238 3836
rect 14238 3780 14294 3836
rect 14294 3780 14298 3836
rect 14234 3776 14298 3780
rect 14314 3836 14378 3840
rect 14314 3780 14318 3836
rect 14318 3780 14374 3836
rect 14374 3780 14378 3836
rect 14314 3776 14378 3780
rect 14394 3836 14458 3840
rect 14394 3780 14398 3836
rect 14398 3780 14454 3836
rect 14454 3780 14458 3836
rect 14394 3776 14458 3780
rect 14474 3836 14538 3840
rect 14474 3780 14478 3836
rect 14478 3780 14534 3836
rect 14534 3780 14538 3836
rect 14474 3776 14538 3780
rect 19547 3836 19611 3840
rect 19547 3780 19551 3836
rect 19551 3780 19607 3836
rect 19607 3780 19611 3836
rect 19547 3776 19611 3780
rect 19627 3836 19691 3840
rect 19627 3780 19631 3836
rect 19631 3780 19687 3836
rect 19687 3780 19691 3836
rect 19627 3776 19691 3780
rect 19707 3836 19771 3840
rect 19707 3780 19711 3836
rect 19711 3780 19767 3836
rect 19767 3780 19771 3836
rect 19707 3776 19771 3780
rect 19787 3836 19851 3840
rect 19787 3780 19791 3836
rect 19791 3780 19847 3836
rect 19847 3780 19851 3836
rect 19787 3776 19851 3780
rect 4268 3292 4332 3296
rect 4268 3236 4272 3292
rect 4272 3236 4328 3292
rect 4328 3236 4332 3292
rect 4268 3232 4332 3236
rect 4348 3292 4412 3296
rect 4348 3236 4352 3292
rect 4352 3236 4408 3292
rect 4408 3236 4412 3292
rect 4348 3232 4412 3236
rect 4428 3292 4492 3296
rect 4428 3236 4432 3292
rect 4432 3236 4488 3292
rect 4488 3236 4492 3292
rect 4428 3232 4492 3236
rect 4508 3292 4572 3296
rect 4508 3236 4512 3292
rect 4512 3236 4568 3292
rect 4568 3236 4572 3292
rect 4508 3232 4572 3236
rect 9581 3292 9645 3296
rect 9581 3236 9585 3292
rect 9585 3236 9641 3292
rect 9641 3236 9645 3292
rect 9581 3232 9645 3236
rect 9661 3292 9725 3296
rect 9661 3236 9665 3292
rect 9665 3236 9721 3292
rect 9721 3236 9725 3292
rect 9661 3232 9725 3236
rect 9741 3292 9805 3296
rect 9741 3236 9745 3292
rect 9745 3236 9801 3292
rect 9801 3236 9805 3292
rect 9741 3232 9805 3236
rect 9821 3292 9885 3296
rect 9821 3236 9825 3292
rect 9825 3236 9881 3292
rect 9881 3236 9885 3292
rect 9821 3232 9885 3236
rect 14894 3292 14958 3296
rect 14894 3236 14898 3292
rect 14898 3236 14954 3292
rect 14954 3236 14958 3292
rect 14894 3232 14958 3236
rect 14974 3292 15038 3296
rect 14974 3236 14978 3292
rect 14978 3236 15034 3292
rect 15034 3236 15038 3292
rect 14974 3232 15038 3236
rect 15054 3292 15118 3296
rect 15054 3236 15058 3292
rect 15058 3236 15114 3292
rect 15114 3236 15118 3292
rect 15054 3232 15118 3236
rect 15134 3292 15198 3296
rect 15134 3236 15138 3292
rect 15138 3236 15194 3292
rect 15194 3236 15198 3292
rect 15134 3232 15198 3236
rect 20207 3292 20271 3296
rect 20207 3236 20211 3292
rect 20211 3236 20267 3292
rect 20267 3236 20271 3292
rect 20207 3232 20271 3236
rect 20287 3292 20351 3296
rect 20287 3236 20291 3292
rect 20291 3236 20347 3292
rect 20347 3236 20351 3292
rect 20287 3232 20351 3236
rect 20367 3292 20431 3296
rect 20367 3236 20371 3292
rect 20371 3236 20427 3292
rect 20427 3236 20431 3292
rect 20367 3232 20431 3236
rect 20447 3292 20511 3296
rect 20447 3236 20451 3292
rect 20451 3236 20507 3292
rect 20507 3236 20511 3292
rect 20447 3232 20511 3236
rect 3608 2748 3672 2752
rect 3608 2692 3612 2748
rect 3612 2692 3668 2748
rect 3668 2692 3672 2748
rect 3608 2688 3672 2692
rect 3688 2748 3752 2752
rect 3688 2692 3692 2748
rect 3692 2692 3748 2748
rect 3748 2692 3752 2748
rect 3688 2688 3752 2692
rect 3768 2748 3832 2752
rect 3768 2692 3772 2748
rect 3772 2692 3828 2748
rect 3828 2692 3832 2748
rect 3768 2688 3832 2692
rect 3848 2748 3912 2752
rect 3848 2692 3852 2748
rect 3852 2692 3908 2748
rect 3908 2692 3912 2748
rect 3848 2688 3912 2692
rect 8921 2748 8985 2752
rect 8921 2692 8925 2748
rect 8925 2692 8981 2748
rect 8981 2692 8985 2748
rect 8921 2688 8985 2692
rect 9001 2748 9065 2752
rect 9001 2692 9005 2748
rect 9005 2692 9061 2748
rect 9061 2692 9065 2748
rect 9001 2688 9065 2692
rect 9081 2748 9145 2752
rect 9081 2692 9085 2748
rect 9085 2692 9141 2748
rect 9141 2692 9145 2748
rect 9081 2688 9145 2692
rect 9161 2748 9225 2752
rect 9161 2692 9165 2748
rect 9165 2692 9221 2748
rect 9221 2692 9225 2748
rect 9161 2688 9225 2692
rect 14234 2748 14298 2752
rect 14234 2692 14238 2748
rect 14238 2692 14294 2748
rect 14294 2692 14298 2748
rect 14234 2688 14298 2692
rect 14314 2748 14378 2752
rect 14314 2692 14318 2748
rect 14318 2692 14374 2748
rect 14374 2692 14378 2748
rect 14314 2688 14378 2692
rect 14394 2748 14458 2752
rect 14394 2692 14398 2748
rect 14398 2692 14454 2748
rect 14454 2692 14458 2748
rect 14394 2688 14458 2692
rect 14474 2748 14538 2752
rect 14474 2692 14478 2748
rect 14478 2692 14534 2748
rect 14534 2692 14538 2748
rect 14474 2688 14538 2692
rect 19547 2748 19611 2752
rect 19547 2692 19551 2748
rect 19551 2692 19607 2748
rect 19607 2692 19611 2748
rect 19547 2688 19611 2692
rect 19627 2748 19691 2752
rect 19627 2692 19631 2748
rect 19631 2692 19687 2748
rect 19687 2692 19691 2748
rect 19627 2688 19691 2692
rect 19707 2748 19771 2752
rect 19707 2692 19711 2748
rect 19711 2692 19767 2748
rect 19767 2692 19771 2748
rect 19707 2688 19771 2692
rect 19787 2748 19851 2752
rect 19787 2692 19791 2748
rect 19791 2692 19847 2748
rect 19847 2692 19851 2748
rect 19787 2688 19851 2692
rect 4268 2204 4332 2208
rect 4268 2148 4272 2204
rect 4272 2148 4328 2204
rect 4328 2148 4332 2204
rect 4268 2144 4332 2148
rect 4348 2204 4412 2208
rect 4348 2148 4352 2204
rect 4352 2148 4408 2204
rect 4408 2148 4412 2204
rect 4348 2144 4412 2148
rect 4428 2204 4492 2208
rect 4428 2148 4432 2204
rect 4432 2148 4488 2204
rect 4488 2148 4492 2204
rect 4428 2144 4492 2148
rect 4508 2204 4572 2208
rect 4508 2148 4512 2204
rect 4512 2148 4568 2204
rect 4568 2148 4572 2204
rect 4508 2144 4572 2148
rect 9581 2204 9645 2208
rect 9581 2148 9585 2204
rect 9585 2148 9641 2204
rect 9641 2148 9645 2204
rect 9581 2144 9645 2148
rect 9661 2204 9725 2208
rect 9661 2148 9665 2204
rect 9665 2148 9721 2204
rect 9721 2148 9725 2204
rect 9661 2144 9725 2148
rect 9741 2204 9805 2208
rect 9741 2148 9745 2204
rect 9745 2148 9801 2204
rect 9801 2148 9805 2204
rect 9741 2144 9805 2148
rect 9821 2204 9885 2208
rect 9821 2148 9825 2204
rect 9825 2148 9881 2204
rect 9881 2148 9885 2204
rect 9821 2144 9885 2148
rect 14894 2204 14958 2208
rect 14894 2148 14898 2204
rect 14898 2148 14954 2204
rect 14954 2148 14958 2204
rect 14894 2144 14958 2148
rect 14974 2204 15038 2208
rect 14974 2148 14978 2204
rect 14978 2148 15034 2204
rect 15034 2148 15038 2204
rect 14974 2144 15038 2148
rect 15054 2204 15118 2208
rect 15054 2148 15058 2204
rect 15058 2148 15114 2204
rect 15114 2148 15118 2204
rect 15054 2144 15118 2148
rect 15134 2204 15198 2208
rect 15134 2148 15138 2204
rect 15138 2148 15194 2204
rect 15194 2148 15198 2204
rect 15134 2144 15198 2148
rect 20207 2204 20271 2208
rect 20207 2148 20211 2204
rect 20211 2148 20267 2204
rect 20267 2148 20271 2204
rect 20207 2144 20271 2148
rect 20287 2204 20351 2208
rect 20287 2148 20291 2204
rect 20291 2148 20347 2204
rect 20347 2148 20351 2204
rect 20287 2144 20351 2148
rect 20367 2204 20431 2208
rect 20367 2148 20371 2204
rect 20371 2148 20427 2204
rect 20427 2148 20431 2204
rect 20367 2144 20431 2148
rect 20447 2204 20511 2208
rect 20447 2148 20451 2204
rect 20451 2148 20507 2204
rect 20507 2148 20511 2204
rect 20447 2144 20511 2148
<< metal4 >>
rect 3600 23424 3920 23440
rect 3600 23360 3608 23424
rect 3672 23360 3688 23424
rect 3752 23360 3768 23424
rect 3832 23360 3848 23424
rect 3912 23360 3920 23424
rect 3600 22336 3920 23360
rect 3600 22272 3608 22336
rect 3672 22272 3688 22336
rect 3752 22272 3768 22336
rect 3832 22272 3848 22336
rect 3912 22272 3920 22336
rect 3600 21248 3920 22272
rect 3600 21184 3608 21248
rect 3672 21184 3688 21248
rect 3752 21184 3768 21248
rect 3832 21184 3848 21248
rect 3912 21184 3920 21248
rect 3600 20858 3920 21184
rect 3600 20622 3642 20858
rect 3878 20622 3920 20858
rect 3600 20160 3920 20622
rect 3600 20096 3608 20160
rect 3672 20096 3688 20160
rect 3752 20096 3768 20160
rect 3832 20096 3848 20160
rect 3912 20096 3920 20160
rect 3600 19072 3920 20096
rect 3600 19008 3608 19072
rect 3672 19008 3688 19072
rect 3752 19008 3768 19072
rect 3832 19008 3848 19072
rect 3912 19008 3920 19072
rect 3600 17984 3920 19008
rect 3600 17920 3608 17984
rect 3672 17920 3688 17984
rect 3752 17920 3768 17984
rect 3832 17920 3848 17984
rect 3912 17920 3920 17984
rect 3600 16896 3920 17920
rect 3600 16832 3608 16896
rect 3672 16832 3688 16896
rect 3752 16832 3768 16896
rect 3832 16832 3848 16896
rect 3912 16832 3920 16896
rect 3600 15808 3920 16832
rect 3600 15744 3608 15808
rect 3672 15744 3688 15808
rect 3752 15744 3768 15808
rect 3832 15744 3848 15808
rect 3912 15744 3920 15808
rect 3600 15554 3920 15744
rect 3600 15318 3642 15554
rect 3878 15318 3920 15554
rect 3600 14720 3920 15318
rect 3600 14656 3608 14720
rect 3672 14656 3688 14720
rect 3752 14656 3768 14720
rect 3832 14656 3848 14720
rect 3912 14656 3920 14720
rect 3600 13632 3920 14656
rect 3600 13568 3608 13632
rect 3672 13568 3688 13632
rect 3752 13568 3768 13632
rect 3832 13568 3848 13632
rect 3912 13568 3920 13632
rect 3600 12544 3920 13568
rect 3600 12480 3608 12544
rect 3672 12480 3688 12544
rect 3752 12480 3768 12544
rect 3832 12480 3848 12544
rect 3912 12480 3920 12544
rect 3600 11456 3920 12480
rect 3600 11392 3608 11456
rect 3672 11392 3688 11456
rect 3752 11392 3768 11456
rect 3832 11392 3848 11456
rect 3912 11392 3920 11456
rect 3600 10368 3920 11392
rect 3600 10304 3608 10368
rect 3672 10304 3688 10368
rect 3752 10304 3768 10368
rect 3832 10304 3848 10368
rect 3912 10304 3920 10368
rect 3600 10250 3920 10304
rect 3600 10014 3642 10250
rect 3878 10014 3920 10250
rect 3600 9280 3920 10014
rect 3600 9216 3608 9280
rect 3672 9216 3688 9280
rect 3752 9216 3768 9280
rect 3832 9216 3848 9280
rect 3912 9216 3920 9280
rect 3600 8192 3920 9216
rect 3600 8128 3608 8192
rect 3672 8128 3688 8192
rect 3752 8128 3768 8192
rect 3832 8128 3848 8192
rect 3912 8128 3920 8192
rect 3600 7104 3920 8128
rect 3600 7040 3608 7104
rect 3672 7040 3688 7104
rect 3752 7040 3768 7104
rect 3832 7040 3848 7104
rect 3912 7040 3920 7104
rect 3600 6016 3920 7040
rect 3600 5952 3608 6016
rect 3672 5952 3688 6016
rect 3752 5952 3768 6016
rect 3832 5952 3848 6016
rect 3912 5952 3920 6016
rect 3600 4946 3920 5952
rect 3600 4928 3642 4946
rect 3878 4928 3920 4946
rect 3600 4864 3608 4928
rect 3912 4864 3920 4928
rect 3600 4710 3642 4864
rect 3878 4710 3920 4864
rect 3600 3840 3920 4710
rect 3600 3776 3608 3840
rect 3672 3776 3688 3840
rect 3752 3776 3768 3840
rect 3832 3776 3848 3840
rect 3912 3776 3920 3840
rect 3600 2752 3920 3776
rect 3600 2688 3608 2752
rect 3672 2688 3688 2752
rect 3752 2688 3768 2752
rect 3832 2688 3848 2752
rect 3912 2688 3920 2752
rect 3600 2128 3920 2688
rect 4260 22880 4580 23440
rect 4260 22816 4268 22880
rect 4332 22816 4348 22880
rect 4412 22816 4428 22880
rect 4492 22816 4508 22880
rect 4572 22816 4580 22880
rect 4260 21792 4580 22816
rect 4260 21728 4268 21792
rect 4332 21728 4348 21792
rect 4412 21728 4428 21792
rect 4492 21728 4508 21792
rect 4572 21728 4580 21792
rect 4260 21518 4580 21728
rect 4260 21282 4302 21518
rect 4538 21282 4580 21518
rect 4260 20704 4580 21282
rect 4260 20640 4268 20704
rect 4332 20640 4348 20704
rect 4412 20640 4428 20704
rect 4492 20640 4508 20704
rect 4572 20640 4580 20704
rect 4260 19616 4580 20640
rect 4260 19552 4268 19616
rect 4332 19552 4348 19616
rect 4412 19552 4428 19616
rect 4492 19552 4508 19616
rect 4572 19552 4580 19616
rect 4260 18528 4580 19552
rect 4260 18464 4268 18528
rect 4332 18464 4348 18528
rect 4412 18464 4428 18528
rect 4492 18464 4508 18528
rect 4572 18464 4580 18528
rect 4260 17440 4580 18464
rect 4260 17376 4268 17440
rect 4332 17376 4348 17440
rect 4412 17376 4428 17440
rect 4492 17376 4508 17440
rect 4572 17376 4580 17440
rect 4260 16352 4580 17376
rect 4260 16288 4268 16352
rect 4332 16288 4348 16352
rect 4412 16288 4428 16352
rect 4492 16288 4508 16352
rect 4572 16288 4580 16352
rect 4260 16214 4580 16288
rect 4260 15978 4302 16214
rect 4538 15978 4580 16214
rect 4260 15264 4580 15978
rect 4260 15200 4268 15264
rect 4332 15200 4348 15264
rect 4412 15200 4428 15264
rect 4492 15200 4508 15264
rect 4572 15200 4580 15264
rect 4260 14176 4580 15200
rect 4260 14112 4268 14176
rect 4332 14112 4348 14176
rect 4412 14112 4428 14176
rect 4492 14112 4508 14176
rect 4572 14112 4580 14176
rect 4260 13088 4580 14112
rect 4260 13024 4268 13088
rect 4332 13024 4348 13088
rect 4412 13024 4428 13088
rect 4492 13024 4508 13088
rect 4572 13024 4580 13088
rect 4260 12000 4580 13024
rect 4260 11936 4268 12000
rect 4332 11936 4348 12000
rect 4412 11936 4428 12000
rect 4492 11936 4508 12000
rect 4572 11936 4580 12000
rect 4260 10912 4580 11936
rect 4260 10848 4268 10912
rect 4332 10910 4348 10912
rect 4412 10910 4428 10912
rect 4492 10910 4508 10912
rect 4572 10848 4580 10912
rect 4260 10674 4302 10848
rect 4538 10674 4580 10848
rect 4260 9824 4580 10674
rect 4260 9760 4268 9824
rect 4332 9760 4348 9824
rect 4412 9760 4428 9824
rect 4492 9760 4508 9824
rect 4572 9760 4580 9824
rect 4260 8736 4580 9760
rect 4260 8672 4268 8736
rect 4332 8672 4348 8736
rect 4412 8672 4428 8736
rect 4492 8672 4508 8736
rect 4572 8672 4580 8736
rect 4260 7648 4580 8672
rect 4260 7584 4268 7648
rect 4332 7584 4348 7648
rect 4412 7584 4428 7648
rect 4492 7584 4508 7648
rect 4572 7584 4580 7648
rect 4260 6560 4580 7584
rect 4260 6496 4268 6560
rect 4332 6496 4348 6560
rect 4412 6496 4428 6560
rect 4492 6496 4508 6560
rect 4572 6496 4580 6560
rect 4260 5606 4580 6496
rect 4260 5472 4302 5606
rect 4538 5472 4580 5606
rect 4260 5408 4268 5472
rect 4572 5408 4580 5472
rect 4260 5370 4302 5408
rect 4538 5370 4580 5408
rect 4260 4384 4580 5370
rect 4260 4320 4268 4384
rect 4332 4320 4348 4384
rect 4412 4320 4428 4384
rect 4492 4320 4508 4384
rect 4572 4320 4580 4384
rect 4260 3296 4580 4320
rect 4260 3232 4268 3296
rect 4332 3232 4348 3296
rect 4412 3232 4428 3296
rect 4492 3232 4508 3296
rect 4572 3232 4580 3296
rect 4260 2208 4580 3232
rect 4260 2144 4268 2208
rect 4332 2144 4348 2208
rect 4412 2144 4428 2208
rect 4492 2144 4508 2208
rect 4572 2144 4580 2208
rect 4260 2128 4580 2144
rect 8913 23424 9233 23440
rect 8913 23360 8921 23424
rect 8985 23360 9001 23424
rect 9065 23360 9081 23424
rect 9145 23360 9161 23424
rect 9225 23360 9233 23424
rect 8913 22336 9233 23360
rect 8913 22272 8921 22336
rect 8985 22272 9001 22336
rect 9065 22272 9081 22336
rect 9145 22272 9161 22336
rect 9225 22272 9233 22336
rect 8913 21248 9233 22272
rect 8913 21184 8921 21248
rect 8985 21184 9001 21248
rect 9065 21184 9081 21248
rect 9145 21184 9161 21248
rect 9225 21184 9233 21248
rect 8913 20858 9233 21184
rect 8913 20622 8955 20858
rect 9191 20622 9233 20858
rect 8913 20160 9233 20622
rect 8913 20096 8921 20160
rect 8985 20096 9001 20160
rect 9065 20096 9081 20160
rect 9145 20096 9161 20160
rect 9225 20096 9233 20160
rect 8913 19072 9233 20096
rect 8913 19008 8921 19072
rect 8985 19008 9001 19072
rect 9065 19008 9081 19072
rect 9145 19008 9161 19072
rect 9225 19008 9233 19072
rect 8913 17984 9233 19008
rect 8913 17920 8921 17984
rect 8985 17920 9001 17984
rect 9065 17920 9081 17984
rect 9145 17920 9161 17984
rect 9225 17920 9233 17984
rect 8913 16896 9233 17920
rect 8913 16832 8921 16896
rect 8985 16832 9001 16896
rect 9065 16832 9081 16896
rect 9145 16832 9161 16896
rect 9225 16832 9233 16896
rect 8913 15808 9233 16832
rect 8913 15744 8921 15808
rect 8985 15744 9001 15808
rect 9065 15744 9081 15808
rect 9145 15744 9161 15808
rect 9225 15744 9233 15808
rect 8913 15554 9233 15744
rect 8913 15318 8955 15554
rect 9191 15318 9233 15554
rect 8913 14720 9233 15318
rect 8913 14656 8921 14720
rect 8985 14656 9001 14720
rect 9065 14656 9081 14720
rect 9145 14656 9161 14720
rect 9225 14656 9233 14720
rect 8913 13632 9233 14656
rect 8913 13568 8921 13632
rect 8985 13568 9001 13632
rect 9065 13568 9081 13632
rect 9145 13568 9161 13632
rect 9225 13568 9233 13632
rect 8913 12544 9233 13568
rect 8913 12480 8921 12544
rect 8985 12480 9001 12544
rect 9065 12480 9081 12544
rect 9145 12480 9161 12544
rect 9225 12480 9233 12544
rect 8913 11456 9233 12480
rect 8913 11392 8921 11456
rect 8985 11392 9001 11456
rect 9065 11392 9081 11456
rect 9145 11392 9161 11456
rect 9225 11392 9233 11456
rect 8913 10368 9233 11392
rect 8913 10304 8921 10368
rect 8985 10304 9001 10368
rect 9065 10304 9081 10368
rect 9145 10304 9161 10368
rect 9225 10304 9233 10368
rect 8913 10250 9233 10304
rect 8913 10014 8955 10250
rect 9191 10014 9233 10250
rect 8913 9280 9233 10014
rect 8913 9216 8921 9280
rect 8985 9216 9001 9280
rect 9065 9216 9081 9280
rect 9145 9216 9161 9280
rect 9225 9216 9233 9280
rect 8913 8192 9233 9216
rect 8913 8128 8921 8192
rect 8985 8128 9001 8192
rect 9065 8128 9081 8192
rect 9145 8128 9161 8192
rect 9225 8128 9233 8192
rect 8913 7104 9233 8128
rect 8913 7040 8921 7104
rect 8985 7040 9001 7104
rect 9065 7040 9081 7104
rect 9145 7040 9161 7104
rect 9225 7040 9233 7104
rect 8913 6016 9233 7040
rect 8913 5952 8921 6016
rect 8985 5952 9001 6016
rect 9065 5952 9081 6016
rect 9145 5952 9161 6016
rect 9225 5952 9233 6016
rect 8913 4946 9233 5952
rect 8913 4928 8955 4946
rect 9191 4928 9233 4946
rect 8913 4864 8921 4928
rect 9225 4864 9233 4928
rect 8913 4710 8955 4864
rect 9191 4710 9233 4864
rect 8913 3840 9233 4710
rect 8913 3776 8921 3840
rect 8985 3776 9001 3840
rect 9065 3776 9081 3840
rect 9145 3776 9161 3840
rect 9225 3776 9233 3840
rect 8913 2752 9233 3776
rect 8913 2688 8921 2752
rect 8985 2688 9001 2752
rect 9065 2688 9081 2752
rect 9145 2688 9161 2752
rect 9225 2688 9233 2752
rect 8913 2128 9233 2688
rect 9573 22880 9893 23440
rect 9573 22816 9581 22880
rect 9645 22816 9661 22880
rect 9725 22816 9741 22880
rect 9805 22816 9821 22880
rect 9885 22816 9893 22880
rect 9573 21792 9893 22816
rect 9573 21728 9581 21792
rect 9645 21728 9661 21792
rect 9725 21728 9741 21792
rect 9805 21728 9821 21792
rect 9885 21728 9893 21792
rect 9573 21518 9893 21728
rect 9573 21282 9615 21518
rect 9851 21282 9893 21518
rect 9573 20704 9893 21282
rect 9573 20640 9581 20704
rect 9645 20640 9661 20704
rect 9725 20640 9741 20704
rect 9805 20640 9821 20704
rect 9885 20640 9893 20704
rect 9573 19616 9893 20640
rect 9573 19552 9581 19616
rect 9645 19552 9661 19616
rect 9725 19552 9741 19616
rect 9805 19552 9821 19616
rect 9885 19552 9893 19616
rect 9573 18528 9893 19552
rect 9573 18464 9581 18528
rect 9645 18464 9661 18528
rect 9725 18464 9741 18528
rect 9805 18464 9821 18528
rect 9885 18464 9893 18528
rect 9573 17440 9893 18464
rect 9573 17376 9581 17440
rect 9645 17376 9661 17440
rect 9725 17376 9741 17440
rect 9805 17376 9821 17440
rect 9885 17376 9893 17440
rect 9573 16352 9893 17376
rect 9573 16288 9581 16352
rect 9645 16288 9661 16352
rect 9725 16288 9741 16352
rect 9805 16288 9821 16352
rect 9885 16288 9893 16352
rect 9573 16214 9893 16288
rect 9573 15978 9615 16214
rect 9851 15978 9893 16214
rect 9573 15264 9893 15978
rect 9573 15200 9581 15264
rect 9645 15200 9661 15264
rect 9725 15200 9741 15264
rect 9805 15200 9821 15264
rect 9885 15200 9893 15264
rect 9573 14176 9893 15200
rect 9573 14112 9581 14176
rect 9645 14112 9661 14176
rect 9725 14112 9741 14176
rect 9805 14112 9821 14176
rect 9885 14112 9893 14176
rect 9573 13088 9893 14112
rect 9573 13024 9581 13088
rect 9645 13024 9661 13088
rect 9725 13024 9741 13088
rect 9805 13024 9821 13088
rect 9885 13024 9893 13088
rect 9573 12000 9893 13024
rect 9573 11936 9581 12000
rect 9645 11936 9661 12000
rect 9725 11936 9741 12000
rect 9805 11936 9821 12000
rect 9885 11936 9893 12000
rect 9573 10912 9893 11936
rect 9573 10848 9581 10912
rect 9645 10910 9661 10912
rect 9725 10910 9741 10912
rect 9805 10910 9821 10912
rect 9885 10848 9893 10912
rect 9573 10674 9615 10848
rect 9851 10674 9893 10848
rect 9573 9824 9893 10674
rect 9573 9760 9581 9824
rect 9645 9760 9661 9824
rect 9725 9760 9741 9824
rect 9805 9760 9821 9824
rect 9885 9760 9893 9824
rect 9573 8736 9893 9760
rect 9573 8672 9581 8736
rect 9645 8672 9661 8736
rect 9725 8672 9741 8736
rect 9805 8672 9821 8736
rect 9885 8672 9893 8736
rect 9573 7648 9893 8672
rect 9573 7584 9581 7648
rect 9645 7584 9661 7648
rect 9725 7584 9741 7648
rect 9805 7584 9821 7648
rect 9885 7584 9893 7648
rect 9573 6560 9893 7584
rect 9573 6496 9581 6560
rect 9645 6496 9661 6560
rect 9725 6496 9741 6560
rect 9805 6496 9821 6560
rect 9885 6496 9893 6560
rect 9573 5606 9893 6496
rect 9573 5472 9615 5606
rect 9851 5472 9893 5606
rect 9573 5408 9581 5472
rect 9885 5408 9893 5472
rect 9573 5370 9615 5408
rect 9851 5370 9893 5408
rect 9573 4384 9893 5370
rect 9573 4320 9581 4384
rect 9645 4320 9661 4384
rect 9725 4320 9741 4384
rect 9805 4320 9821 4384
rect 9885 4320 9893 4384
rect 9573 3296 9893 4320
rect 9573 3232 9581 3296
rect 9645 3232 9661 3296
rect 9725 3232 9741 3296
rect 9805 3232 9821 3296
rect 9885 3232 9893 3296
rect 9573 2208 9893 3232
rect 9573 2144 9581 2208
rect 9645 2144 9661 2208
rect 9725 2144 9741 2208
rect 9805 2144 9821 2208
rect 9885 2144 9893 2208
rect 9573 2128 9893 2144
rect 14226 23424 14546 23440
rect 14226 23360 14234 23424
rect 14298 23360 14314 23424
rect 14378 23360 14394 23424
rect 14458 23360 14474 23424
rect 14538 23360 14546 23424
rect 14226 22336 14546 23360
rect 14226 22272 14234 22336
rect 14298 22272 14314 22336
rect 14378 22272 14394 22336
rect 14458 22272 14474 22336
rect 14538 22272 14546 22336
rect 14226 21248 14546 22272
rect 14226 21184 14234 21248
rect 14298 21184 14314 21248
rect 14378 21184 14394 21248
rect 14458 21184 14474 21248
rect 14538 21184 14546 21248
rect 14226 20858 14546 21184
rect 14226 20622 14268 20858
rect 14504 20622 14546 20858
rect 14226 20160 14546 20622
rect 14226 20096 14234 20160
rect 14298 20096 14314 20160
rect 14378 20096 14394 20160
rect 14458 20096 14474 20160
rect 14538 20096 14546 20160
rect 14226 19072 14546 20096
rect 14226 19008 14234 19072
rect 14298 19008 14314 19072
rect 14378 19008 14394 19072
rect 14458 19008 14474 19072
rect 14538 19008 14546 19072
rect 14226 17984 14546 19008
rect 14226 17920 14234 17984
rect 14298 17920 14314 17984
rect 14378 17920 14394 17984
rect 14458 17920 14474 17984
rect 14538 17920 14546 17984
rect 14226 16896 14546 17920
rect 14226 16832 14234 16896
rect 14298 16832 14314 16896
rect 14378 16832 14394 16896
rect 14458 16832 14474 16896
rect 14538 16832 14546 16896
rect 14226 15808 14546 16832
rect 14226 15744 14234 15808
rect 14298 15744 14314 15808
rect 14378 15744 14394 15808
rect 14458 15744 14474 15808
rect 14538 15744 14546 15808
rect 14226 15554 14546 15744
rect 14226 15318 14268 15554
rect 14504 15318 14546 15554
rect 14226 14720 14546 15318
rect 14226 14656 14234 14720
rect 14298 14656 14314 14720
rect 14378 14656 14394 14720
rect 14458 14656 14474 14720
rect 14538 14656 14546 14720
rect 14226 13632 14546 14656
rect 14226 13568 14234 13632
rect 14298 13568 14314 13632
rect 14378 13568 14394 13632
rect 14458 13568 14474 13632
rect 14538 13568 14546 13632
rect 14226 12544 14546 13568
rect 14226 12480 14234 12544
rect 14298 12480 14314 12544
rect 14378 12480 14394 12544
rect 14458 12480 14474 12544
rect 14538 12480 14546 12544
rect 14226 11456 14546 12480
rect 14226 11392 14234 11456
rect 14298 11392 14314 11456
rect 14378 11392 14394 11456
rect 14458 11392 14474 11456
rect 14538 11392 14546 11456
rect 14226 10368 14546 11392
rect 14226 10304 14234 10368
rect 14298 10304 14314 10368
rect 14378 10304 14394 10368
rect 14458 10304 14474 10368
rect 14538 10304 14546 10368
rect 14226 10250 14546 10304
rect 14226 10014 14268 10250
rect 14504 10014 14546 10250
rect 14226 9280 14546 10014
rect 14226 9216 14234 9280
rect 14298 9216 14314 9280
rect 14378 9216 14394 9280
rect 14458 9216 14474 9280
rect 14538 9216 14546 9280
rect 14226 8192 14546 9216
rect 14226 8128 14234 8192
rect 14298 8128 14314 8192
rect 14378 8128 14394 8192
rect 14458 8128 14474 8192
rect 14538 8128 14546 8192
rect 14226 7104 14546 8128
rect 14226 7040 14234 7104
rect 14298 7040 14314 7104
rect 14378 7040 14394 7104
rect 14458 7040 14474 7104
rect 14538 7040 14546 7104
rect 14226 6016 14546 7040
rect 14226 5952 14234 6016
rect 14298 5952 14314 6016
rect 14378 5952 14394 6016
rect 14458 5952 14474 6016
rect 14538 5952 14546 6016
rect 14226 4946 14546 5952
rect 14226 4928 14268 4946
rect 14504 4928 14546 4946
rect 14226 4864 14234 4928
rect 14538 4864 14546 4928
rect 14226 4710 14268 4864
rect 14504 4710 14546 4864
rect 14226 3840 14546 4710
rect 14226 3776 14234 3840
rect 14298 3776 14314 3840
rect 14378 3776 14394 3840
rect 14458 3776 14474 3840
rect 14538 3776 14546 3840
rect 14226 2752 14546 3776
rect 14226 2688 14234 2752
rect 14298 2688 14314 2752
rect 14378 2688 14394 2752
rect 14458 2688 14474 2752
rect 14538 2688 14546 2752
rect 14226 2128 14546 2688
rect 14886 22880 15206 23440
rect 14886 22816 14894 22880
rect 14958 22816 14974 22880
rect 15038 22816 15054 22880
rect 15118 22816 15134 22880
rect 15198 22816 15206 22880
rect 14886 21792 15206 22816
rect 14886 21728 14894 21792
rect 14958 21728 14974 21792
rect 15038 21728 15054 21792
rect 15118 21728 15134 21792
rect 15198 21728 15206 21792
rect 14886 21518 15206 21728
rect 14886 21282 14928 21518
rect 15164 21282 15206 21518
rect 14886 20704 15206 21282
rect 14886 20640 14894 20704
rect 14958 20640 14974 20704
rect 15038 20640 15054 20704
rect 15118 20640 15134 20704
rect 15198 20640 15206 20704
rect 14886 19616 15206 20640
rect 14886 19552 14894 19616
rect 14958 19552 14974 19616
rect 15038 19552 15054 19616
rect 15118 19552 15134 19616
rect 15198 19552 15206 19616
rect 14886 18528 15206 19552
rect 14886 18464 14894 18528
rect 14958 18464 14974 18528
rect 15038 18464 15054 18528
rect 15118 18464 15134 18528
rect 15198 18464 15206 18528
rect 14886 17440 15206 18464
rect 14886 17376 14894 17440
rect 14958 17376 14974 17440
rect 15038 17376 15054 17440
rect 15118 17376 15134 17440
rect 15198 17376 15206 17440
rect 14886 16352 15206 17376
rect 14886 16288 14894 16352
rect 14958 16288 14974 16352
rect 15038 16288 15054 16352
rect 15118 16288 15134 16352
rect 15198 16288 15206 16352
rect 14886 16214 15206 16288
rect 14886 15978 14928 16214
rect 15164 15978 15206 16214
rect 14886 15264 15206 15978
rect 14886 15200 14894 15264
rect 14958 15200 14974 15264
rect 15038 15200 15054 15264
rect 15118 15200 15134 15264
rect 15198 15200 15206 15264
rect 14886 14176 15206 15200
rect 14886 14112 14894 14176
rect 14958 14112 14974 14176
rect 15038 14112 15054 14176
rect 15118 14112 15134 14176
rect 15198 14112 15206 14176
rect 14886 13088 15206 14112
rect 14886 13024 14894 13088
rect 14958 13024 14974 13088
rect 15038 13024 15054 13088
rect 15118 13024 15134 13088
rect 15198 13024 15206 13088
rect 14886 12000 15206 13024
rect 14886 11936 14894 12000
rect 14958 11936 14974 12000
rect 15038 11936 15054 12000
rect 15118 11936 15134 12000
rect 15198 11936 15206 12000
rect 14886 10912 15206 11936
rect 14886 10848 14894 10912
rect 14958 10910 14974 10912
rect 15038 10910 15054 10912
rect 15118 10910 15134 10912
rect 15198 10848 15206 10912
rect 14886 10674 14928 10848
rect 15164 10674 15206 10848
rect 14886 9824 15206 10674
rect 14886 9760 14894 9824
rect 14958 9760 14974 9824
rect 15038 9760 15054 9824
rect 15118 9760 15134 9824
rect 15198 9760 15206 9824
rect 14886 8736 15206 9760
rect 14886 8672 14894 8736
rect 14958 8672 14974 8736
rect 15038 8672 15054 8736
rect 15118 8672 15134 8736
rect 15198 8672 15206 8736
rect 14886 7648 15206 8672
rect 14886 7584 14894 7648
rect 14958 7584 14974 7648
rect 15038 7584 15054 7648
rect 15118 7584 15134 7648
rect 15198 7584 15206 7648
rect 14886 6560 15206 7584
rect 14886 6496 14894 6560
rect 14958 6496 14974 6560
rect 15038 6496 15054 6560
rect 15118 6496 15134 6560
rect 15198 6496 15206 6560
rect 14886 5606 15206 6496
rect 14886 5472 14928 5606
rect 15164 5472 15206 5606
rect 14886 5408 14894 5472
rect 15198 5408 15206 5472
rect 14886 5370 14928 5408
rect 15164 5370 15206 5408
rect 14886 4384 15206 5370
rect 14886 4320 14894 4384
rect 14958 4320 14974 4384
rect 15038 4320 15054 4384
rect 15118 4320 15134 4384
rect 15198 4320 15206 4384
rect 14886 3296 15206 4320
rect 14886 3232 14894 3296
rect 14958 3232 14974 3296
rect 15038 3232 15054 3296
rect 15118 3232 15134 3296
rect 15198 3232 15206 3296
rect 14886 2208 15206 3232
rect 14886 2144 14894 2208
rect 14958 2144 14974 2208
rect 15038 2144 15054 2208
rect 15118 2144 15134 2208
rect 15198 2144 15206 2208
rect 14886 2128 15206 2144
rect 19539 23424 19859 23440
rect 19539 23360 19547 23424
rect 19611 23360 19627 23424
rect 19691 23360 19707 23424
rect 19771 23360 19787 23424
rect 19851 23360 19859 23424
rect 19539 22336 19859 23360
rect 19539 22272 19547 22336
rect 19611 22272 19627 22336
rect 19691 22272 19707 22336
rect 19771 22272 19787 22336
rect 19851 22272 19859 22336
rect 19539 21248 19859 22272
rect 19539 21184 19547 21248
rect 19611 21184 19627 21248
rect 19691 21184 19707 21248
rect 19771 21184 19787 21248
rect 19851 21184 19859 21248
rect 19539 20858 19859 21184
rect 19539 20622 19581 20858
rect 19817 20622 19859 20858
rect 19539 20160 19859 20622
rect 19539 20096 19547 20160
rect 19611 20096 19627 20160
rect 19691 20096 19707 20160
rect 19771 20096 19787 20160
rect 19851 20096 19859 20160
rect 19539 19072 19859 20096
rect 19539 19008 19547 19072
rect 19611 19008 19627 19072
rect 19691 19008 19707 19072
rect 19771 19008 19787 19072
rect 19851 19008 19859 19072
rect 19539 17984 19859 19008
rect 19539 17920 19547 17984
rect 19611 17920 19627 17984
rect 19691 17920 19707 17984
rect 19771 17920 19787 17984
rect 19851 17920 19859 17984
rect 19539 16896 19859 17920
rect 19539 16832 19547 16896
rect 19611 16832 19627 16896
rect 19691 16832 19707 16896
rect 19771 16832 19787 16896
rect 19851 16832 19859 16896
rect 19539 15808 19859 16832
rect 19539 15744 19547 15808
rect 19611 15744 19627 15808
rect 19691 15744 19707 15808
rect 19771 15744 19787 15808
rect 19851 15744 19859 15808
rect 19539 15554 19859 15744
rect 19539 15318 19581 15554
rect 19817 15318 19859 15554
rect 19539 14720 19859 15318
rect 19539 14656 19547 14720
rect 19611 14656 19627 14720
rect 19691 14656 19707 14720
rect 19771 14656 19787 14720
rect 19851 14656 19859 14720
rect 19539 13632 19859 14656
rect 19539 13568 19547 13632
rect 19611 13568 19627 13632
rect 19691 13568 19707 13632
rect 19771 13568 19787 13632
rect 19851 13568 19859 13632
rect 19539 12544 19859 13568
rect 19539 12480 19547 12544
rect 19611 12480 19627 12544
rect 19691 12480 19707 12544
rect 19771 12480 19787 12544
rect 19851 12480 19859 12544
rect 19539 11456 19859 12480
rect 19539 11392 19547 11456
rect 19611 11392 19627 11456
rect 19691 11392 19707 11456
rect 19771 11392 19787 11456
rect 19851 11392 19859 11456
rect 19539 10368 19859 11392
rect 19539 10304 19547 10368
rect 19611 10304 19627 10368
rect 19691 10304 19707 10368
rect 19771 10304 19787 10368
rect 19851 10304 19859 10368
rect 19539 10250 19859 10304
rect 19539 10014 19581 10250
rect 19817 10014 19859 10250
rect 19539 9280 19859 10014
rect 19539 9216 19547 9280
rect 19611 9216 19627 9280
rect 19691 9216 19707 9280
rect 19771 9216 19787 9280
rect 19851 9216 19859 9280
rect 19539 8192 19859 9216
rect 19539 8128 19547 8192
rect 19611 8128 19627 8192
rect 19691 8128 19707 8192
rect 19771 8128 19787 8192
rect 19851 8128 19859 8192
rect 19539 7104 19859 8128
rect 19539 7040 19547 7104
rect 19611 7040 19627 7104
rect 19691 7040 19707 7104
rect 19771 7040 19787 7104
rect 19851 7040 19859 7104
rect 19539 6016 19859 7040
rect 19539 5952 19547 6016
rect 19611 5952 19627 6016
rect 19691 5952 19707 6016
rect 19771 5952 19787 6016
rect 19851 5952 19859 6016
rect 19539 4946 19859 5952
rect 19539 4928 19581 4946
rect 19817 4928 19859 4946
rect 19539 4864 19547 4928
rect 19851 4864 19859 4928
rect 19539 4710 19581 4864
rect 19817 4710 19859 4864
rect 19539 3840 19859 4710
rect 19539 3776 19547 3840
rect 19611 3776 19627 3840
rect 19691 3776 19707 3840
rect 19771 3776 19787 3840
rect 19851 3776 19859 3840
rect 19539 2752 19859 3776
rect 19539 2688 19547 2752
rect 19611 2688 19627 2752
rect 19691 2688 19707 2752
rect 19771 2688 19787 2752
rect 19851 2688 19859 2752
rect 19539 2128 19859 2688
rect 20199 22880 20519 23440
rect 20199 22816 20207 22880
rect 20271 22816 20287 22880
rect 20351 22816 20367 22880
rect 20431 22816 20447 22880
rect 20511 22816 20519 22880
rect 20199 21792 20519 22816
rect 20199 21728 20207 21792
rect 20271 21728 20287 21792
rect 20351 21728 20367 21792
rect 20431 21728 20447 21792
rect 20511 21728 20519 21792
rect 20199 21518 20519 21728
rect 20199 21282 20241 21518
rect 20477 21282 20519 21518
rect 20199 20704 20519 21282
rect 20199 20640 20207 20704
rect 20271 20640 20287 20704
rect 20351 20640 20367 20704
rect 20431 20640 20447 20704
rect 20511 20640 20519 20704
rect 20199 19616 20519 20640
rect 20199 19552 20207 19616
rect 20271 19552 20287 19616
rect 20351 19552 20367 19616
rect 20431 19552 20447 19616
rect 20511 19552 20519 19616
rect 20199 18528 20519 19552
rect 20199 18464 20207 18528
rect 20271 18464 20287 18528
rect 20351 18464 20367 18528
rect 20431 18464 20447 18528
rect 20511 18464 20519 18528
rect 20199 17440 20519 18464
rect 20199 17376 20207 17440
rect 20271 17376 20287 17440
rect 20351 17376 20367 17440
rect 20431 17376 20447 17440
rect 20511 17376 20519 17440
rect 20199 16352 20519 17376
rect 20199 16288 20207 16352
rect 20271 16288 20287 16352
rect 20351 16288 20367 16352
rect 20431 16288 20447 16352
rect 20511 16288 20519 16352
rect 20199 16214 20519 16288
rect 20199 15978 20241 16214
rect 20477 15978 20519 16214
rect 20199 15264 20519 15978
rect 20199 15200 20207 15264
rect 20271 15200 20287 15264
rect 20351 15200 20367 15264
rect 20431 15200 20447 15264
rect 20511 15200 20519 15264
rect 20199 14176 20519 15200
rect 20199 14112 20207 14176
rect 20271 14112 20287 14176
rect 20351 14112 20367 14176
rect 20431 14112 20447 14176
rect 20511 14112 20519 14176
rect 20199 13088 20519 14112
rect 20199 13024 20207 13088
rect 20271 13024 20287 13088
rect 20351 13024 20367 13088
rect 20431 13024 20447 13088
rect 20511 13024 20519 13088
rect 20199 12000 20519 13024
rect 20199 11936 20207 12000
rect 20271 11936 20287 12000
rect 20351 11936 20367 12000
rect 20431 11936 20447 12000
rect 20511 11936 20519 12000
rect 20199 10912 20519 11936
rect 20199 10848 20207 10912
rect 20271 10910 20287 10912
rect 20351 10910 20367 10912
rect 20431 10910 20447 10912
rect 20511 10848 20519 10912
rect 20199 10674 20241 10848
rect 20477 10674 20519 10848
rect 20199 9824 20519 10674
rect 20199 9760 20207 9824
rect 20271 9760 20287 9824
rect 20351 9760 20367 9824
rect 20431 9760 20447 9824
rect 20511 9760 20519 9824
rect 20199 8736 20519 9760
rect 20199 8672 20207 8736
rect 20271 8672 20287 8736
rect 20351 8672 20367 8736
rect 20431 8672 20447 8736
rect 20511 8672 20519 8736
rect 20199 7648 20519 8672
rect 20199 7584 20207 7648
rect 20271 7584 20287 7648
rect 20351 7584 20367 7648
rect 20431 7584 20447 7648
rect 20511 7584 20519 7648
rect 20199 6560 20519 7584
rect 20199 6496 20207 6560
rect 20271 6496 20287 6560
rect 20351 6496 20367 6560
rect 20431 6496 20447 6560
rect 20511 6496 20519 6560
rect 20199 5606 20519 6496
rect 20199 5472 20241 5606
rect 20477 5472 20519 5606
rect 20199 5408 20207 5472
rect 20511 5408 20519 5472
rect 20199 5370 20241 5408
rect 20477 5370 20519 5408
rect 20199 4384 20519 5370
rect 20199 4320 20207 4384
rect 20271 4320 20287 4384
rect 20351 4320 20367 4384
rect 20431 4320 20447 4384
rect 20511 4320 20519 4384
rect 20199 3296 20519 4320
rect 20199 3232 20207 3296
rect 20271 3232 20287 3296
rect 20351 3232 20367 3296
rect 20431 3232 20447 3296
rect 20511 3232 20519 3296
rect 20199 2208 20519 3232
rect 20199 2144 20207 2208
rect 20271 2144 20287 2208
rect 20351 2144 20367 2208
rect 20431 2144 20447 2208
rect 20511 2144 20519 2208
rect 20199 2128 20519 2144
<< via4 >>
rect 3642 20622 3878 20858
rect 3642 15318 3878 15554
rect 3642 10014 3878 10250
rect 3642 4928 3878 4946
rect 3642 4864 3672 4928
rect 3672 4864 3688 4928
rect 3688 4864 3752 4928
rect 3752 4864 3768 4928
rect 3768 4864 3832 4928
rect 3832 4864 3848 4928
rect 3848 4864 3878 4928
rect 3642 4710 3878 4864
rect 4302 21282 4538 21518
rect 4302 15978 4538 16214
rect 4302 10848 4332 10910
rect 4332 10848 4348 10910
rect 4348 10848 4412 10910
rect 4412 10848 4428 10910
rect 4428 10848 4492 10910
rect 4492 10848 4508 10910
rect 4508 10848 4538 10910
rect 4302 10674 4538 10848
rect 4302 5472 4538 5606
rect 4302 5408 4332 5472
rect 4332 5408 4348 5472
rect 4348 5408 4412 5472
rect 4412 5408 4428 5472
rect 4428 5408 4492 5472
rect 4492 5408 4508 5472
rect 4508 5408 4538 5472
rect 4302 5370 4538 5408
rect 8955 20622 9191 20858
rect 8955 15318 9191 15554
rect 8955 10014 9191 10250
rect 8955 4928 9191 4946
rect 8955 4864 8985 4928
rect 8985 4864 9001 4928
rect 9001 4864 9065 4928
rect 9065 4864 9081 4928
rect 9081 4864 9145 4928
rect 9145 4864 9161 4928
rect 9161 4864 9191 4928
rect 8955 4710 9191 4864
rect 9615 21282 9851 21518
rect 9615 15978 9851 16214
rect 9615 10848 9645 10910
rect 9645 10848 9661 10910
rect 9661 10848 9725 10910
rect 9725 10848 9741 10910
rect 9741 10848 9805 10910
rect 9805 10848 9821 10910
rect 9821 10848 9851 10910
rect 9615 10674 9851 10848
rect 9615 5472 9851 5606
rect 9615 5408 9645 5472
rect 9645 5408 9661 5472
rect 9661 5408 9725 5472
rect 9725 5408 9741 5472
rect 9741 5408 9805 5472
rect 9805 5408 9821 5472
rect 9821 5408 9851 5472
rect 9615 5370 9851 5408
rect 14268 20622 14504 20858
rect 14268 15318 14504 15554
rect 14268 10014 14504 10250
rect 14268 4928 14504 4946
rect 14268 4864 14298 4928
rect 14298 4864 14314 4928
rect 14314 4864 14378 4928
rect 14378 4864 14394 4928
rect 14394 4864 14458 4928
rect 14458 4864 14474 4928
rect 14474 4864 14504 4928
rect 14268 4710 14504 4864
rect 14928 21282 15164 21518
rect 14928 15978 15164 16214
rect 14928 10848 14958 10910
rect 14958 10848 14974 10910
rect 14974 10848 15038 10910
rect 15038 10848 15054 10910
rect 15054 10848 15118 10910
rect 15118 10848 15134 10910
rect 15134 10848 15164 10910
rect 14928 10674 15164 10848
rect 14928 5472 15164 5606
rect 14928 5408 14958 5472
rect 14958 5408 14974 5472
rect 14974 5408 15038 5472
rect 15038 5408 15054 5472
rect 15054 5408 15118 5472
rect 15118 5408 15134 5472
rect 15134 5408 15164 5472
rect 14928 5370 15164 5408
rect 19581 20622 19817 20858
rect 19581 15318 19817 15554
rect 19581 10014 19817 10250
rect 19581 4928 19817 4946
rect 19581 4864 19611 4928
rect 19611 4864 19627 4928
rect 19627 4864 19691 4928
rect 19691 4864 19707 4928
rect 19707 4864 19771 4928
rect 19771 4864 19787 4928
rect 19787 4864 19817 4928
rect 19581 4710 19817 4864
rect 20241 21282 20477 21518
rect 20241 15978 20477 16214
rect 20241 10848 20271 10910
rect 20271 10848 20287 10910
rect 20287 10848 20351 10910
rect 20351 10848 20367 10910
rect 20367 10848 20431 10910
rect 20431 10848 20447 10910
rect 20447 10848 20477 10910
rect 20241 10674 20477 10848
rect 20241 5472 20477 5606
rect 20241 5408 20271 5472
rect 20271 5408 20287 5472
rect 20287 5408 20351 5472
rect 20351 5408 20367 5472
rect 20367 5408 20431 5472
rect 20431 5408 20447 5472
rect 20447 5408 20477 5472
rect 20241 5370 20477 5408
<< metal5 >>
rect 1056 21518 22404 21560
rect 1056 21282 4302 21518
rect 4538 21282 9615 21518
rect 9851 21282 14928 21518
rect 15164 21282 20241 21518
rect 20477 21282 22404 21518
rect 1056 21240 22404 21282
rect 1056 20858 22404 20900
rect 1056 20622 3642 20858
rect 3878 20622 8955 20858
rect 9191 20622 14268 20858
rect 14504 20622 19581 20858
rect 19817 20622 22404 20858
rect 1056 20580 22404 20622
rect 1056 16214 22404 16256
rect 1056 15978 4302 16214
rect 4538 15978 9615 16214
rect 9851 15978 14928 16214
rect 15164 15978 20241 16214
rect 20477 15978 22404 16214
rect 1056 15936 22404 15978
rect 1056 15554 22404 15596
rect 1056 15318 3642 15554
rect 3878 15318 8955 15554
rect 9191 15318 14268 15554
rect 14504 15318 19581 15554
rect 19817 15318 22404 15554
rect 1056 15276 22404 15318
rect 1056 10910 22404 10952
rect 1056 10674 4302 10910
rect 4538 10674 9615 10910
rect 9851 10674 14928 10910
rect 15164 10674 20241 10910
rect 20477 10674 22404 10910
rect 1056 10632 22404 10674
rect 1056 10250 22404 10292
rect 1056 10014 3642 10250
rect 3878 10014 8955 10250
rect 9191 10014 14268 10250
rect 14504 10014 19581 10250
rect 19817 10014 22404 10250
rect 1056 9972 22404 10014
rect 1056 5606 22404 5648
rect 1056 5370 4302 5606
rect 4538 5370 9615 5606
rect 9851 5370 14928 5606
rect 15164 5370 20241 5606
rect 20477 5370 22404 5606
rect 1056 5328 22404 5370
rect 1056 4946 22404 4988
rect 1056 4710 3642 4946
rect 3878 4710 8955 4946
rect 9191 4710 14268 4946
rect 14504 4710 19581 4946
rect 19817 4710 22404 4946
rect 1056 4668 22404 4710
use sky130_fd_sc_hd__nor4_1  _1388_
timestamp 0
transform 1 0 15364 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _1389_
timestamp 0
transform -1 0 18216 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__nor4_1  _1390_
timestamp 0
transform -1 0 8280 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1391_
timestamp 0
transform -1 0 7728 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _1392_
timestamp 0
transform 1 0 12328 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1393_
timestamp 0
transform 1 0 13616 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1394_
timestamp 0
transform -1 0 15456 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_4  _1395_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__nor4_1  _1396_
timestamp 0
transform -1 0 6808 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _1397_
timestamp 0
transform -1 0 13248 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1398_
timestamp 0
transform -1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1399_
timestamp 0
transform 1 0 13248 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  _1400_
timestamp 0
transform -1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1401_
timestamp 0
transform 1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1402_
timestamp 0
transform -1 0 8832 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1403_
timestamp 0
transform -1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1404_
timestamp 0
transform 1 0 9936 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1405_
timestamp 0
transform 1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _1406_
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_0  _1407_
timestamp 0
transform 1 0 11776 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1408_
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _1409_
timestamp 0
transform -1 0 11684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _1410_
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _1411_
timestamp 0
transform -1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _1412_
timestamp 0
transform -1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1413_
timestamp 0
transform -1 0 9660 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1414_
timestamp 0
transform -1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1415_
timestamp 0
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1416_
timestamp 0
transform 1 0 12788 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1417_
timestamp 0
transform 1 0 12328 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1418_
timestamp 0
transform 1 0 12972 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1419_
timestamp 0
transform -1 0 12144 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1420_
timestamp 0
transform 1 0 12144 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1421_
timestamp 0
transform 1 0 12788 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1422_
timestamp 0
transform -1 0 13248 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1423_
timestamp 0
transform 1 0 11868 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1424_
timestamp 0
transform -1 0 12512 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1425__150
timestamp 0
transform -1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _1425_
timestamp 0
transform -1 0 13800 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _1426_
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1427_
timestamp 0
transform 1 0 12604 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1428_
timestamp 0
transform -1 0 3588 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1429_
timestamp 0
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1430_
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1431_
timestamp 0
transform 1 0 2392 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1432_
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1433_
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1434_
timestamp 0
transform 1 0 2944 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1435_
timestamp 0
transform -1 0 5060 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1436_
timestamp 0
transform 1 0 5060 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1437_
timestamp 0
transform -1 0 3312 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1438_
timestamp 0
transform -1 0 2484 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1439__151
timestamp 0
transform -1 0 5888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1439_
timestamp 0
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1440_
timestamp 0
transform -1 0 5980 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1441_
timestamp 0
transform -1 0 4600 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1442_
timestamp 0
transform -1 0 2760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1443_
timestamp 0
transform 1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1444_
timestamp 0
transform 1 0 4232 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1445_
timestamp 0
transform 1 0 2392 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1446_
timestamp 0
transform 1 0 4692 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1447_
timestamp 0
transform 1 0 2852 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1448_
timestamp 0
transform 1 0 2760 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1449_
timestamp 0
transform 1 0 3772 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1450_
timestamp 0
transform 1 0 3864 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1451_
timestamp 0
transform -1 0 2944 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1452_
timestamp 0
transform -1 0 2484 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1453__152
timestamp 0
transform -1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1453_
timestamp 0
transform -1 0 5612 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1454_
timestamp 0
transform -1 0 6440 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1455_
timestamp 0
transform -1 0 3772 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1456_
timestamp 0
transform -1 0 5888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1457_
timestamp 0
transform -1 0 4600 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1458_
timestamp 0
transform 1 0 5612 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1459_
timestamp 0
transform -1 0 5888 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1460_
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1461_
timestamp 0
transform 1 0 3864 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1462_
timestamp 0
transform 1 0 4324 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1463_
timestamp 0
transform 1 0 4968 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1464_
timestamp 0
transform 1 0 4968 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1465_
timestamp 0
transform 1 0 4784 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1466_
timestamp 0
transform 1 0 4048 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1467__153
timestamp 0
transform -1 0 6992 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 0
transform 1 0 5520 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1468_
timestamp 0
transform -1 0 6164 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1469_
timestamp 0
transform -1 0 5796 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1470_
timestamp 0
transform -1 0 8464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1471_
timestamp 0
transform -1 0 8740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1472_
timestamp 0
transform -1 0 8648 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1473_
timestamp 0
transform 1 0 6900 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1474_
timestamp 0
transform -1 0 8372 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1475_
timestamp 0
transform 1 0 8372 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1476_
timestamp 0
transform 1 0 6900 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1477_
timestamp 0
transform 1 0 7268 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1478_
timestamp 0
transform 1 0 7084 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1479_
timestamp 0
transform 1 0 7544 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1480_
timestamp 0
transform 1 0 7360 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1481__154
timestamp 0
transform -1 0 8280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1481_
timestamp 0
transform 1 0 7176 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1482_
timestamp 0
transform -1 0 7820 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1483_
timestamp 0
transform 1 0 7360 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1484_
timestamp 0
transform -1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1485_
timestamp 0
transform -1 0 11776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1486_
timestamp 0
transform -1 0 10488 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1487_
timestamp 0
transform 1 0 11500 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1488_
timestamp 0
transform 1 0 10580 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1489_
timestamp 0
transform -1 0 9752 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1490_
timestamp 0
transform -1 0 10304 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1491_
timestamp 0
transform 1 0 9292 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1492_
timestamp 0
transform -1 0 9568 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 0
transform 1 0 10672 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1494_
timestamp 0
transform 1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1495__155
timestamp 0
transform 1 0 8096 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1495_
timestamp 0
transform 1 0 8372 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1496_
timestamp 0
transform 1 0 7912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1497_
timestamp 0
transform 1 0 9752 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1498_
timestamp 0
transform -1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1499_
timestamp 0
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1500_
timestamp 0
transform -1 0 10764 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1501_
timestamp 0
transform 1 0 10764 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1502_
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1503_
timestamp 0
transform 1 0 10672 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1504_
timestamp 0
transform -1 0 10672 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1505_
timestamp 0
transform 1 0 10488 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1506_
timestamp 0
transform -1 0 10488 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 0
transform 1 0 10580 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 0
transform 1 0 10488 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1509__156
timestamp 0
transform -1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1509_
timestamp 0
transform 1 0 8464 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1510_
timestamp 0
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1511_
timestamp 0
transform 1 0 9476 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1512_
timestamp 0
transform -1 0 13616 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1513_
timestamp 0
transform -1 0 13248 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1514_
timestamp 0
transform 1 0 13064 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1515_
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1516_
timestamp 0
transform 1 0 13156 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1517_
timestamp 0
transform 1 0 12696 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1518_
timestamp 0
transform 1 0 12604 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1519_
timestamp 0
transform -1 0 12604 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1520_
timestamp 0
transform 1 0 13248 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 0
transform 1 0 13064 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 0
transform -1 0 13064 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1523__157
timestamp 0
transform -1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 0
transform 1 0 14996 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 0
transform -1 0 15640 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 0
transform -1 0 14352 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1526_
timestamp 0
transform -1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1527_
timestamp 0
transform -1 0 13800 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1528_
timestamp 0
transform 1 0 13524 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1529_
timestamp 0
transform -1 0 12696 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1530_
timestamp 0
transform 1 0 13432 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1531_
timestamp 0
transform 1 0 13248 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1532_
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1533_
timestamp 0
transform 1 0 13064 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1534_
timestamp 0
transform 1 0 12880 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1535_
timestamp 0
transform 1 0 12696 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1536_
timestamp 0
transform 1 0 12604 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1537__158
timestamp 0
transform -1 0 13984 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1537_
timestamp 0
transform 1 0 12880 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1538_
timestamp 0
transform -1 0 12880 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1539_
timestamp 0
transform 1 0 12696 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1540_
timestamp 0
transform 1 0 15180 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1541_
timestamp 0
transform -1 0 16560 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1542_
timestamp 0
transform -1 0 14996 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1543_
timestamp 0
transform -1 0 16376 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1544_
timestamp 0
transform 1 0 15916 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1545_
timestamp 0
transform 1 0 15456 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1546_
timestamp 0
transform -1 0 16468 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1547_
timestamp 0
transform 1 0 15180 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1548_
timestamp 0
transform -1 0 15548 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1549_
timestamp 0
transform 1 0 15640 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1550_
timestamp 0
transform 1 0 15456 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1551__128
timestamp 0
transform -1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 0
transform 1 0 14812 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1552_
timestamp 0
transform 1 0 14260 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 0
transform 1 0 14996 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1554_
timestamp 0
transform -1 0 20332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1555_
timestamp 0
transform -1 0 20332 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1556_
timestamp 0
transform -1 0 18676 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1557_
timestamp 0
transform -1 0 19136 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1558_
timestamp 0
transform -1 0 18952 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1559_
timestamp 0
transform -1 0 19228 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1560_
timestamp 0
transform -1 0 18492 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1561_
timestamp 0
transform 1 0 17388 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1562_
timestamp 0
transform -1 0 17388 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1563_
timestamp 0
transform 1 0 19228 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1564_
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1565__129
timestamp 0
transform -1 0 17480 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1565_
timestamp 0
transform -1 0 17204 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1566_
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 0
transform 1 0 17940 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1568_
timestamp 0
transform 1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1569_
timestamp 0
transform -1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1570_
timestamp 0
transform -1 0 10580 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1571_
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1572_
timestamp 0
transform 1 0 9568 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1573_
timestamp 0
transform -1 0 9476 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1574_
timestamp 0
transform -1 0 10948 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1575_
timestamp 0
transform 1 0 10396 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1576_
timestamp 0
transform -1 0 10396 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1577_
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1578_
timestamp 0
transform 1 0 9384 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1579__130
timestamp 0
transform -1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1579_
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1580_
timestamp 0
transform 1 0 8832 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1581_
timestamp 0
transform 1 0 9476 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1582_
timestamp 0
transform -1 0 21252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1583_
timestamp 0
transform -1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1584_
timestamp 0
transform -1 0 19780 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1585_
timestamp 0
transform -1 0 19964 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1586_
timestamp 0
transform -1 0 19136 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1587_
timestamp 0
transform -1 0 19320 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1588_
timestamp 0
transform -1 0 19872 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1589_
timestamp 0
transform 1 0 18400 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1590_
timestamp 0
transform -1 0 18676 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1591_
timestamp 0
transform 1 0 20148 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1592_
timestamp 0
transform 1 0 19964 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1593__131
timestamp 0
transform 1 0 17940 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1593_
timestamp 0
transform 1 0 17664 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1594_
timestamp 0
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1595_
timestamp 0
transform 1 0 18676 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1596_
timestamp 0
transform 1 0 20424 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1597_
timestamp 0
transform -1 0 20608 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1598_
timestamp 0
transform -1 0 19688 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1599_
timestamp 0
transform -1 0 18308 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1600_
timestamp 0
transform -1 0 18952 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1601_
timestamp 0
transform -1 0 19044 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1602_
timestamp 0
transform -1 0 19780 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1603_
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1604_
timestamp 0
transform -1 0 19044 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1605_
timestamp 0
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1606_
timestamp 0
transform 1 0 19872 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1607__132
timestamp 0
transform -1 0 19136 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1607_
timestamp 0
transform 1 0 18032 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1608_
timestamp 0
transform 1 0 17204 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1609_
timestamp 0
transform 1 0 18308 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1610_
timestamp 0
transform -1 0 17756 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1611_
timestamp 0
transform -1 0 16376 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1612_
timestamp 0
transform 1 0 17480 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1613_
timestamp 0
transform -1 0 17480 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1614_
timestamp 0
transform 1 0 16100 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1615_
timestamp 0
transform 1 0 15180 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1616_
timestamp 0
transform 1 0 14904 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1617_
timestamp 0
transform -1 0 16100 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1618_
timestamp 0
transform 1 0 15732 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1619_
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1620_
timestamp 0
transform 1 0 15272 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1621__133
timestamp 0
transform -1 0 16468 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 0
transform 1 0 15732 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1622_
timestamp 0
transform 1 0 15272 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1623_
timestamp 0
transform 1 0 15548 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1624_
timestamp 0
transform -1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1625_
timestamp 0
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1626_
timestamp 0
transform -1 0 11776 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1627_
timestamp 0
transform 1 0 11776 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1628_
timestamp 0
transform 1 0 13616 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1629_
timestamp 0
transform 1 0 13064 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1630_
timestamp 0
transform 1 0 12604 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1631_
timestamp 0
transform -1 0 13984 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1632_
timestamp 0
transform -1 0 13984 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1633_
timestamp 0
transform -1 0 13064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1634_
timestamp 0
transform -1 0 12604 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1635__134
timestamp 0
transform -1 0 13708 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1635_
timestamp 0
transform 1 0 13064 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1636_
timestamp 0
transform -1 0 13064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1637_
timestamp 0
transform -1 0 13064 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1638_
timestamp 0
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1639_
timestamp 0
transform 1 0 13248 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1640_
timestamp 0
transform 1 0 13800 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1641_
timestamp 0
transform 1 0 14904 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1642_
timestamp 0
transform 1 0 15824 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1643_
timestamp 0
transform 1 0 13524 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1644_
timestamp 0
transform 1 0 14076 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1645_
timestamp 0
transform 1 0 15364 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1646_
timestamp 0
transform 1 0 14260 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 0
transform 1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1648_
timestamp 0
transform -1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1649__135
timestamp 0
transform 1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1649_
timestamp 0
transform 1 0 15088 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 0
transform -1 0 15088 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1651_
timestamp 0
transform -1 0 15088 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1652_
timestamp 0
transform 1 0 19688 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1653_
timestamp 0
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1654_
timestamp 0
transform -1 0 18952 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1655_
timestamp 0
transform -1 0 18768 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1656_
timestamp 0
transform 1 0 18676 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1657_
timestamp 0
transform 1 0 18032 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1658_
timestamp 0
transform -1 0 18032 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1659_
timestamp 0
transform 1 0 18216 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1660_
timestamp 0
transform 1 0 17572 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1661_
timestamp 0
transform 1 0 20056 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1662_
timestamp 0
transform 1 0 19228 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1663__136
timestamp 0
transform 1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1663_
timestamp 0
transform 1 0 17480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1664_
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 0
transform 1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1666_
timestamp 0
transform 1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1667_
timestamp 0
transform -1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1668_
timestamp 0
transform 1 0 20240 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1669_
timestamp 0
transform 1 0 19228 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1670_
timestamp 0
transform -1 0 20240 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1671_
timestamp 0
transform 1 0 19688 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1672_
timestamp 0
transform -1 0 19780 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1673_
timestamp 0
transform 1 0 18400 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1674_
timestamp 0
transform -1 0 19136 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 0
transform 1 0 20884 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1676_
timestamp 0
transform 1 0 20056 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1677__137
timestamp 0
transform -1 0 18492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 0
transform 1 0 17664 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 0
transform 1 0 16836 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1680_
timestamp 0
transform -1 0 21620 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1681_
timestamp 0
transform -1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1682_
timestamp 0
transform -1 0 19228 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1683_
timestamp 0
transform -1 0 20332 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1684_
timestamp 0
transform -1 0 18768 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1685_
timestamp 0
transform -1 0 20332 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1686_
timestamp 0
transform -1 0 19872 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1687_
timestamp 0
transform -1 0 19412 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1688_
timestamp 0
transform -1 0 19136 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 0
transform 1 0 20424 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 0
transform 1 0 20240 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1691__138
timestamp 0
transform 1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1691_
timestamp 0
transform 1 0 17204 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1692_
timestamp 0
transform 1 0 16376 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1693_
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1694_
timestamp 0
transform -1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1695_
timestamp 0
transform -1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1696_
timestamp 0
transform -1 0 18124 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1697_
timestamp 0
transform -1 0 19688 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1698_
timestamp 0
transform 1 0 18584 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1699_
timestamp 0
transform 1 0 18124 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1700_
timestamp 0
transform -1 0 19688 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1701_
timestamp 0
transform -1 0 19136 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1702_
timestamp 0
transform -1 0 19044 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 0
transform 1 0 19964 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1704_
timestamp 0
transform 1 0 18768 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1705__139
timestamp 0
transform -1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 0
transform 1 0 17664 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1706_
timestamp 0
transform 1 0 16836 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1707_
timestamp 0
transform 1 0 18216 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1708_
timestamp 0
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1709_
timestamp 0
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1710_
timestamp 0
transform 1 0 16652 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1711_
timestamp 0
transform -1 0 15916 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1712_
timestamp 0
transform 1 0 16928 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1713_
timestamp 0
transform 1 0 16192 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1714_
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1715_
timestamp 0
transform -1 0 16928 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1716_
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 0
transform 1 0 17480 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1718_
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1719_
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1719__140
timestamp 0
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1720_
timestamp 0
transform 1 0 15548 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1721_
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1722_
timestamp 0
transform -1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1723_
timestamp 0
transform 1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1724_
timestamp 0
transform 1 0 6992 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1725_
timestamp 0
transform 1 0 6992 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1726_
timestamp 0
transform 1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1727_
timestamp 0
transform -1 0 6256 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1728_
timestamp 0
transform 1 0 6440 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1729_
timestamp 0
transform 1 0 8004 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1730_
timestamp 0
transform 1 0 7360 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1731_
timestamp 0
transform 1 0 7084 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1732_
timestamp 0
transform 1 0 6624 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1733__141
timestamp 0
transform -1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 0
transform 1 0 7544 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1734_
timestamp 0
transform -1 0 8096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1735_
timestamp 0
transform -1 0 7912 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1736_
timestamp 0
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1737_
timestamp 0
transform -1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1738_
timestamp 0
transform 1 0 13064 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1739_
timestamp 0
transform 1 0 13524 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1740_
timestamp 0
transform 1 0 13524 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1741_
timestamp 0
transform 1 0 12880 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1742_
timestamp 0
transform 1 0 13340 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1743_
timestamp 0
transform -1 0 14536 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1744_
timestamp 0
transform -1 0 15732 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1745_
timestamp 0
transform 1 0 14628 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 0
transform 1 0 13800 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1747__142
timestamp 0
transform -1 0 15180 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1747_
timestamp 0
transform 1 0 14444 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1748_
timestamp 0
transform 1 0 14076 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1749_
timestamp 0
transform -1 0 14812 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1750_
timestamp 0
transform -1 0 6256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1751_
timestamp 0
transform 1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1752_
timestamp 0
transform 1 0 3864 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1753_
timestamp 0
transform 1 0 4324 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1754_
timestamp 0
transform 1 0 4048 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1755_
timestamp 0
transform -1 0 3680 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1756_
timestamp 0
transform 1 0 4600 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1757_
timestamp 0
transform -1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1758_
timestamp 0
transform 1 0 5520 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 0
transform 1 0 4048 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1760_
timestamp 0
transform -1 0 4600 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1761__143
timestamp 0
transform 1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1762_
timestamp 0
transform -1 0 6624 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 0
transform -1 0 5336 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1764_
timestamp 0
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1765_
timestamp 0
transform -1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1766_
timestamp 0
transform 1 0 3220 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1767_
timestamp 0
transform 1 0 2760 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1768_
timestamp 0
transform 1 0 4048 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1769_
timestamp 0
transform 1 0 3128 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1770_
timestamp 0
transform 1 0 3036 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1771_
timestamp 0
transform -1 0 5060 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1772_
timestamp 0
transform 1 0 4600 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 0
transform -1 0 3128 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1774_
timestamp 0
transform -1 0 2300 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1775__144
timestamp 0
transform -1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 0
transform -1 0 5888 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 0
transform -1 0 4600 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1778_
timestamp 0
transform -1 0 3036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1779_
timestamp 0
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1780_
timestamp 0
transform -1 0 2024 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1781_
timestamp 0
transform 1 0 2852 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1782_
timestamp 0
transform 1 0 4508 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1783_
timestamp 0
transform 1 0 3036 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1784_
timestamp 0
transform 1 0 3680 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1785_
timestamp 0
transform 1 0 4232 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1786_
timestamp 0
transform 1 0 3956 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 0
transform -1 0 2852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1788_
timestamp 0
transform -1 0 2760 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1789__145
timestamp 0
transform -1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1790_
timestamp 0
transform -1 0 5428 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1791_
timestamp 0
transform -1 0 3680 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1792_
timestamp 0
transform -1 0 8096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1793_
timestamp 0
transform -1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1794_
timestamp 0
transform 1 0 6532 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1795_
timestamp 0
transform 1 0 8004 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1796_
timestamp 0
transform 1 0 7636 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1797_
timestamp 0
transform -1 0 8004 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1798_
timestamp 0
transform 1 0 6624 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1799_
timestamp 0
transform 1 0 7360 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1800_
timestamp 0
transform 1 0 6716 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 0
transform 1 0 6992 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 0
transform 1 0 6900 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1803__146
timestamp 0
transform 1 0 6716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1803_
timestamp 0
transform 1 0 6808 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 0
transform -1 0 6808 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1805_
timestamp 0
transform 1 0 6716 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1806_
timestamp 0
transform -1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1807_
timestamp 0
transform 1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1808_
timestamp 0
transform -1 0 10948 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1809_
timestamp 0
transform 1 0 10396 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1810_
timestamp 0
transform -1 0 9844 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1811_
timestamp 0
transform -1 0 10396 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1812_
timestamp 0
transform -1 0 10488 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1813_
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1814_
timestamp 0
transform 1 0 9016 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1815_
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1816_
timestamp 0
transform 1 0 11960 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1817__147
timestamp 0
transform -1 0 10120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 0
transform 1 0 9016 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1818_
timestamp 0
transform 1 0 8740 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 0
transform 1 0 10212 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1820_
timestamp 0
transform -1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1821_
timestamp 0
transform -1 0 11224 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1822_
timestamp 0
transform -1 0 9844 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1823_
timestamp 0
transform -1 0 9384 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1824_
timestamp 0
transform 1 0 9384 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1825_
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1826_
timestamp 0
transform 1 0 8924 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1827_
timestamp 0
transform 1 0 9844 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1828_
timestamp 0
transform -1 0 8924 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1829_
timestamp 0
transform 1 0 9844 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1830_
timestamp 0
transform 1 0 9844 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1831__148
timestamp 0
transform -1 0 8832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1831_
timestamp 0
transform 1 0 7728 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1832_
timestamp 0
transform 1 0 7728 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1833_
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1834_
timestamp 0
transform 1 0 4600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1835_
timestamp 0
transform -1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1836_
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1837_
timestamp 0
transform -1 0 5980 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1838_
timestamp 0
transform -1 0 4876 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1839_
timestamp 0
transform -1 0 5612 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1840_
timestamp 0
transform 1 0 4048 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1841_
timestamp 0
transform -1 0 6072 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1842_
timestamp 0
transform -1 0 6992 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1843_
timestamp 0
transform -1 0 5152 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1844_
timestamp 0
transform -1 0 4324 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1845__149
timestamp 0
transform -1 0 7268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1845_
timestamp 0
transform 1 0 6164 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1846_
timestamp 0
transform -1 0 6164 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1847_
timestamp 0
transform -1 0 5520 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1910_
timestamp 0
transform 1 0 7636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1911_
timestamp 0
transform -1 0 8648 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1912_
timestamp 0
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1913_
timestamp 0
transform 1 0 6440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1914_
timestamp 0
transform -1 0 7452 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1915_
timestamp 0
transform 1 0 5428 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1916_
timestamp 0
transform 1 0 6440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1917_
timestamp 0
transform 1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1918_
timestamp 0
transform 1 0 7544 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1919_
timestamp 0
transform 1 0 6256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1920_
timestamp 0
transform 1 0 6808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1921_
timestamp 0
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1922_
timestamp 0
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1923_
timestamp 0
transform 1 0 7176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1924_
timestamp 0
transform -1 0 7820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1925_
timestamp 0
transform 1 0 6992 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1926_
timestamp 0
transform -1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1927_
timestamp 0
transform 1 0 13524 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1928_
timestamp 0
transform -1 0 14076 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1929_
timestamp 0
transform -1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1930_
timestamp 0
transform -1 0 16376 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1931_
timestamp 0
transform -1 0 16560 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1932_
timestamp 0
transform -1 0 16100 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1933_
timestamp 0
transform 1 0 12420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1934_
timestamp 0
transform -1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1935_
timestamp 0
transform -1 0 16744 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1936_
timestamp 0
transform -1 0 16560 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1937_
timestamp 0
transform -1 0 15916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1938_
timestamp 0
transform -1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1939_
timestamp 0
transform -1 0 15364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1940_
timestamp 0
transform -1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1941_
timestamp 0
transform -1 0 16192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clone1
timestamp 0
transform -1 0 11408 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clone2
timestamp 0
transform 1 0 6992 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout107
timestamp 0
transform -1 0 6072 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 0
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout109
timestamp 0
transform 1 0 4784 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 0
transform -1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout111
timestamp 0
transform 1 0 5336 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout112
timestamp 0
transform -1 0 3680 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout113
timestamp 0
transform 1 0 15732 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp 0
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout115
timestamp 0
transform 1 0 4876 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout116
timestamp 0
transform -1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout117
timestamp 0
transform 1 0 12512 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 0
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout119
timestamp 0
transform 1 0 4968 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout120
timestamp 0
transform -1 0 2852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  fanout121
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout122
timestamp 0
transform 1 0 4876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout123
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  fanout124
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout125
timestamp 0
transform -1 0 14904 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout126
timestamp 0
transform -1 0 3404 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout127
timestamp 0
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_23
timestamp 0
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_34
timestamp 0
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_48
timestamp 0
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77
timestamp 0
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_90
timestamp 0
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_104
timestamp 0
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_118
timestamp 0
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_135
timestamp 0
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 0
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_147
timestamp 0
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_161
timestamp 0
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_175
timestamp 0
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_188
timestamp 0
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_202
timestamp 0
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 0
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_77
timestamp 0
transform 1 0 8188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_89
timestamp 0
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_97
timestamp 0
transform 1 0 10028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 0
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_133
timestamp 0
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_156
timestamp 0
transform 1 0 15456 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_164
timestamp 0
transform 1 0 16192 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_187
timestamp 0
transform 1 0 18308 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_199
timestamp 0
transform 1 0 19412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_211
timestamp 0
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_7
timestamp 0
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 0
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_49
timestamp 0
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_56
timestamp 0
transform 1 0 6256 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_69
timestamp 0
transform 1 0 7452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 0
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_89
timestamp 0
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_99
timestamp 0
transform 1 0 10212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_114
timestamp 0
transform 1 0 11592 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_126
timestamp 0
transform 1 0 12696 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_150
timestamp 0
transform 1 0 14904 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_162
timestamp 0
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_200
timestamp 0
transform 1 0 19504 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_212
timestamp 0
transform 1 0 20608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_224
timestamp 0
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_31
timestamp 0
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_74
timestamp 0
transform 1 0 7912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_86
timestamp 0
transform 1 0 9016 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_92
timestamp 0
transform 1 0 9568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_103
timestamp 0
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_122
timestamp 0
transform 1 0 12328 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_155
timestamp 0
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_178
timestamp 0
transform 1 0 17480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_190
timestamp 0
transform 1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_201
timestamp 0
transform 1 0 19596 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_213
timestamp 0
transform 1 0 20700 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_221
timestamp 0
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 0
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 0
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 0
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_59
timestamp 0
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_63
timestamp 0
transform 1 0 6900 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_69
timestamp 0
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 0
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_107
timestamp 0
transform 1 0 10948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_119
timestamp 0
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_131
timestamp 0
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_165
timestamp 0
transform 1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_177
timestamp 0
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 0
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_202
timestamp 0
transform 1 0 19688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_217
timestamp 0
transform 1 0 21068 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 0
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_40
timestamp 0
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_49
timestamp 0
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_61
timestamp 0
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_67
timestamp 0
transform 1 0 7268 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_80
timestamp 0
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_97
timestamp 0
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 0
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_124
timestamp 0
transform 1 0 12512 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_136
timestamp 0
transform 1 0 13616 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_146
timestamp 0
transform 1 0 14536 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_158
timestamp 0
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 0
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_183
timestamp 0
transform 1 0 17940 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_202
timestamp 0
transform 1 0 19688 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_214
timestamp 0
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 0
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_7
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_19
timestamp 0
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_45
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_55
timestamp 0
transform 1 0 6164 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_67
timestamp 0
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_79
timestamp 0
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_93
timestamp 0
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_108
timestamp 0
transform 1 0 11040 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_134
timestamp 0
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_154
timestamp 0
transform 1 0 15272 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_166
timestamp 0
transform 1 0 16376 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_178
timestamp 0
transform 1 0 17480 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_190
timestamp 0
transform 1 0 18584 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 0
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_221
timestamp 0
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_6
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_18
timestamp 0
transform 1 0 2760 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_26
timestamp 0
transform 1 0 3496 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_31
timestamp 0
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_52
timestamp 0
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_66
timestamp 0
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_79
timestamp 0
transform 1 0 8372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_83
timestamp 0
transform 1 0 8740 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_139
timestamp 0
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_153
timestamp 0
transform 1 0 15180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_178
timestamp 0
transform 1 0 17480 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_186
timestamp 0
transform 1 0 18216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_195
timestamp 0
transform 1 0 19044 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_203
timestamp 0
transform 1 0 19780 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_209
timestamp 0
transform 1 0 20332 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_217
timestamp 0
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_48
timestamp 0
transform 1 0 5520 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_63
timestamp 0
transform 1 0 6900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_75
timestamp 0
transform 1 0 8004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 0
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_132
timestamp 0
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_166
timestamp 0
transform 1 0 16376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_170
timestamp 0
transform 1 0 16744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_192
timestamp 0
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_209
timestamp 0
transform 1 0 20332 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_219
timestamp 0
transform 1 0 21252 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_227
timestamp 0
transform 1 0 21988 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 0
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_13
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_19
timestamp 0
transform 1 0 2852 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_28
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 0
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_74
timestamp 0
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_86
timestamp 0
transform 1 0 9016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_94
timestamp 0
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_101
timestamp 0
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 0
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_121
timestamp 0
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_132
timestamp 0
transform 1 0 13248 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_144
timestamp 0
transform 1 0 14352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_148
timestamp 0
transform 1 0 14720 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_155
timestamp 0
transform 1 0 15364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_204
timestamp 0
transform 1 0 19872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 0
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_38
timestamp 0
transform 1 0 4600 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_57
timestamp 0
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_61
timestamp 0
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_69
timestamp 0
transform 1 0 7452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_78
timestamp 0
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 0
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_145
timestamp 0
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_156
timestamp 0
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_161
timestamp 0
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_165
timestamp 0
transform 1 0 16284 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_184
timestamp 0
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_188
timestamp 0
transform 1 0 18400 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_206
timestamp 0
transform 1 0 20056 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_218
timestamp 0
transform 1 0 21160 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_7
timestamp 0
transform 1 0 1748 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_28
timestamp 0
transform 1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_37
timestamp 0
transform 1 0 4508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_45
timestamp 0
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 0
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_78
timestamp 0
transform 1 0 8280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 0
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_138
timestamp 0
transform 1 0 13800 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_146
timestamp 0
transform 1 0 14536 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_150
timestamp 0
transform 1 0 14904 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_162
timestamp 0
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_172
timestamp 0
transform 1 0 16928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_176
timestamp 0
transform 1 0 17296 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_180
timestamp 0
transform 1 0 17664 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_192
timestamp 0
transform 1 0 18768 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_206
timestamp 0
transform 1 0 20056 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_218
timestamp 0
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_225
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_7
timestamp 0
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_19
timestamp 0
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_74
timestamp 0
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 0
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_118
timestamp 0
transform 1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 0
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_164
timestamp 0
transform 1 0 16192 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_176
timestamp 0
transform 1 0 17296 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 0
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 0
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_221
timestamp 0
transform 1 0 21436 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_33
timestamp 0
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 0
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 0
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_74
timestamp 0
transform 1 0 7912 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_86
timestamp 0
transform 1 0 9016 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_98
timestamp 0
transform 1 0 10120 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 0
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_149
timestamp 0
transform 1 0 14812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_157
timestamp 0
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_216
timestamp 0
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_7
timestamp 0
transform 1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 0
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_50
timestamp 0
transform 1 0 5704 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_106
timestamp 0
transform 1 0 10856 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_118
timestamp 0
transform 1 0 11960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_132
timestamp 0
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_152
timestamp 0
transform 1 0 15088 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_164
timestamp 0
transform 1 0 16192 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_170
timestamp 0
transform 1 0 16744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_35
timestamp 0
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 0
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_75
timestamp 0
transform 1 0 8004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_120
timestamp 0
transform 1 0 12144 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_132
timestamp 0
transform 1 0 13248 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_155
timestamp 0
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_193
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_207
timestamp 0
transform 1 0 20148 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_212
timestamp 0
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_42
timestamp 0
transform 1 0 4968 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_46
timestamp 0
transform 1 0 5336 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_58
timestamp 0
transform 1 0 6440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_67
timestamp 0
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_76
timestamp 0
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_98
timestamp 0
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_108
timestamp 0
transform 1 0 11040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_127
timestamp 0
transform 1 0 12788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_131
timestamp 0
transform 1 0 13156 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_162
timestamp 0
transform 1 0 16008 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_170
timestamp 0
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 0
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_221
timestamp 0
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_9
timestamp 0
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_13
timestamp 0
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_25
timestamp 0
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_37
timestamp 0
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_49
timestamp 0
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_80
timestamp 0
transform 1 0 8464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_107
timestamp 0
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_117
timestamp 0
transform 1 0 11868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_129
timestamp 0
transform 1 0 12972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 0
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_192
timestamp 0
transform 1 0 18768 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_204
timestamp 0
transform 1 0 19872 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_216
timestamp 0
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_33
timestamp 0
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 0
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp 0
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_89
timestamp 0
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_95
timestamp 0
transform 1 0 9844 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_101
timestamp 0
transform 1 0 10396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_113
timestamp 0
transform 1 0 11500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_127
timestamp 0
transform 1 0 12788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_165
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_176
timestamp 0
transform 1 0 17296 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 0
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_197
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_205
timestamp 0
transform 1 0 19964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_217
timestamp 0
transform 1 0 21068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_225
timestamp 0
transform 1 0 21804 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_6
timestamp 0
transform 1 0 1656 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_18
timestamp 0
transform 1 0 2760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_49
timestamp 0
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_75
timestamp 0
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_87
timestamp 0
transform 1 0 9108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_99
timestamp 0
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_117
timestamp 0
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_135
timestamp 0
transform 1 0 13524 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_141
timestamp 0
transform 1 0 14076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_153
timestamp 0
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 0
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_181
timestamp 0
transform 1 0 17756 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_194
timestamp 0
transform 1 0 18952 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_215
timestamp 0
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 0
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_6
timestamp 0
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_18
timestamp 0
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 0
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_58
timestamp 0
transform 1 0 6440 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_70
timestamp 0
transform 1 0 7544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 0
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_104
timestamp 0
transform 1 0 10672 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_110
timestamp 0
transform 1 0 11224 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_132
timestamp 0
transform 1 0 13248 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_166
timestamp 0
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_178
timestamp 0
transform 1 0 17480 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_190
timestamp 0
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 0
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_221
timestamp 0
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_6
timestamp 0
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 0
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_30
timestamp 0
transform 1 0 3864 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 0
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_64
timestamp 0
transform 1 0 6992 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_76
timestamp 0
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_92
timestamp 0
transform 1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 0
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_130
timestamp 0
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_140
timestamp 0
transform 1 0 13984 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_152
timestamp 0
transform 1 0 15088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 0
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_195
timestamp 0
transform 1 0 19044 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_207
timestamp 0
transform 1 0 20148 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_219
timestamp 0
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 0
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_6
timestamp 0
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_18
timestamp 0
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 0
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_45
timestamp 0
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_67
timestamp 0
transform 1 0 7268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_79
timestamp 0
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_102
timestamp 0
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_114
timestamp 0
transform 1 0 11592 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_122
timestamp 0
transform 1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_148
timestamp 0
transform 1 0 14720 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_183
timestamp 0
transform 1 0 17940 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 0
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_202
timestamp 0
transform 1 0 19688 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_208
timestamp 0
transform 1 0 20240 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_212
timestamp 0
transform 1 0 20608 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_224
timestamp 0
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_12
timestamp 0
transform 1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_32
timestamp 0
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_50
timestamp 0
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_90
timestamp 0
transform 1 0 9384 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_102
timestamp 0
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 0
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_130
timestamp 0
transform 1 0 13064 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_157
timestamp 0
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 0
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_203
timestamp 0
transform 1 0 19780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 0
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_225
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_38
timestamp 0
transform 1 0 4600 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_59
timestamp 0
transform 1 0 6532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_71
timestamp 0
transform 1 0 7636 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_101
timestamp 0
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_111
timestamp 0
transform 1 0 11316 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_126
timestamp 0
transform 1 0 12696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 0
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_168
timestamp 0
transform 1 0 16560 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_180
timestamp 0
transform 1 0 17664 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_204
timestamp 0
transform 1 0 19872 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_213
timestamp 0
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_7
timestamp 0
transform 1 0 1748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_13
timestamp 0
transform 1 0 2300 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_25
timestamp 0
transform 1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_32
timestamp 0
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_44
timestamp 0
transform 1 0 5152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 0
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_65
timestamp 0
transform 1 0 7084 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_77
timestamp 0
transform 1 0 8188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_85
timestamp 0
transform 1 0 8924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_97
timestamp 0
transform 1 0 10028 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_116
timestamp 0
transform 1 0 11776 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_128
timestamp 0
transform 1 0 12880 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_132
timestamp 0
transform 1 0 13248 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_136
timestamp 0
transform 1 0 13616 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_148
timestamp 0
transform 1 0 14720 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_163
timestamp 0
transform 1 0 16100 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_196
timestamp 0
transform 1 0 19136 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_208
timestamp 0
transform 1 0 20240 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_220
timestamp 0
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_6
timestamp 0
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_18
timestamp 0
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 0
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_52
timestamp 0
transform 1 0 5888 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_67
timestamp 0
transform 1 0 7268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 0
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_110
timestamp 0
transform 1 0 11224 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_118
timestamp 0
transform 1 0 11960 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_163
timestamp 0
transform 1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_168
timestamp 0
transform 1 0 16560 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_180
timestamp 0
transform 1 0 17664 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_192
timestamp 0
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_221
timestamp 0
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_7
timestamp 0
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_19
timestamp 0
transform 1 0 2852 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_31
timestamp 0
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_43
timestamp 0
transform 1 0 5060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_51
timestamp 0
transform 1 0 5796 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_77
timestamp 0
transform 1 0 8188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_89
timestamp 0
transform 1 0 9292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 0
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_144
timestamp 0
transform 1 0 14352 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_148
timestamp 0
transform 1 0 14720 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_187
timestamp 0
transform 1 0 18308 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_203
timestamp 0
transform 1 0 19780 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_215
timestamp 0
transform 1 0 20884 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_219
timestamp 0
transform 1 0 21252 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_25
timestamp 0
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_37
timestamp 0
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_58
timestamp 0
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_62
timestamp 0
transform 1 0 6808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_66
timestamp 0
transform 1 0 7176 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_72
timestamp 0
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_88
timestamp 0
transform 1 0 9200 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_94
timestamp 0
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_114
timestamp 0
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_149
timestamp 0
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_163
timestamp 0
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_175
timestamp 0
transform 1 0 17204 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_183
timestamp 0
transform 1 0 17940 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_204
timestamp 0
transform 1 0 19872 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_219
timestamp 0
transform 1 0 21252 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_227
timestamp 0
transform 1 0 21988 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_7
timestamp 0
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_36
timestamp 0
transform 1 0 4416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_65
timestamp 0
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_73
timestamp 0
transform 1 0 7820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_85
timestamp 0
transform 1 0 8924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_97
timestamp 0
transform 1 0 10028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 0
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_141
timestamp 0
transform 1 0 14076 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_153
timestamp 0
transform 1 0 15180 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_159
timestamp 0
transform 1 0 15732 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 0
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_189
timestamp 0
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_217
timestamp 0
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_6
timestamp 0
transform 1 0 1656 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_24
timestamp 0
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_33
timestamp 0
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_47
timestamp 0
transform 1 0 5428 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_64
timestamp 0
transform 1 0 6992 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_72
timestamp 0
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_102
timestamp 0
transform 1 0 10488 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_114
timestamp 0
transform 1 0 11592 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_126
timestamp 0
transform 1 0 12696 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 0
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 0
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_177
timestamp 0
transform 1 0 17388 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_186
timestamp 0
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 0
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 0
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_221
timestamp 0
transform 1 0 21436 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_7
timestamp 0
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_19
timestamp 0
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_31
timestamp 0
transform 1 0 3956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_39
timestamp 0
transform 1 0 4692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_49
timestamp 0
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 0
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_63
timestamp 0
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_73
timestamp 0
transform 1 0 7820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_88
timestamp 0
transform 1 0 9200 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_108
timestamp 0
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_116
timestamp 0
transform 1 0 11776 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_141
timestamp 0
transform 1 0 14076 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_152
timestamp 0
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_164
timestamp 0
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_178
timestamp 0
transform 1 0 17480 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_190
timestamp 0
transform 1 0 18584 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_202
timestamp 0
transform 1 0 19688 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_214
timestamp 0
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 0
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 0
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 0
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_41
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_54
timestamp 0
transform 1 0 6072 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_78
timestamp 0
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_92
timestamp 0
transform 1 0 9568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_100
timestamp 0
transform 1 0 10304 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_118
timestamp 0
transform 1 0 11960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_178
timestamp 0
transform 1 0 17480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 0
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 0
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_221
timestamp 0
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_72
timestamp 0
transform 1 0 7728 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_84
timestamp 0
transform 1 0 8832 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_88
timestamp 0
transform 1 0 9200 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_96
timestamp 0
transform 1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_100
timestamp 0
transform 1 0 10304 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 0
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_116
timestamp 0
transform 1 0 11776 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_128
timestamp 0
transform 1 0 12880 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 0
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_149
timestamp 0
transform 1 0 14812 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_157
timestamp 0
transform 1 0 15548 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 0
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_177
timestamp 0
transform 1 0 17388 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_209
timestamp 0
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 0
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_7
timestamp 0
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 0
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_52
timestamp 0
transform 1 0 5888 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_64
timestamp 0
transform 1 0 6992 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_72
timestamp 0
transform 1 0 7728 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_79
timestamp 0
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 0
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_133
timestamp 0
transform 1 0 13340 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_158
timestamp 0
transform 1 0 15640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_166
timestamp 0
transform 1 0 16376 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_174
timestamp 0
transform 1 0 17112 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_184
timestamp 0
transform 1 0 18032 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_221
timestamp 0
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_7
timestamp 0
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_19
timestamp 0
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_31
timestamp 0
transform 1 0 3956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_38
timestamp 0
transform 1 0 4600 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_52
timestamp 0
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_84
timestamp 0
transform 1 0 8832 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_96
timestamp 0
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_108
timestamp 0
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_155
timestamp 0
transform 1 0 15364 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 0
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 0
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 0
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 0
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 0
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_6
timestamp 0
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_18
timestamp 0
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 0
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_61
timestamp 0
transform 1 0 6716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_82
timestamp 0
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 0
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_144
timestamp 0
transform 1 0 14352 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_167
timestamp 0
transform 1 0 16468 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_179
timestamp 0
transform 1 0 17572 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_191
timestamp 0
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_221
timestamp 0
transform 1 0 21436 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_227
timestamp 0
transform 1 0 21988 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_12
timestamp 0
transform 1 0 2208 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_24
timestamp 0
transform 1 0 3312 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_36
timestamp 0
transform 1 0 4416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_48
timestamp 0
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_65
timestamp 0
transform 1 0 7084 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_83
timestamp 0
transform 1 0 8740 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_95
timestamp 0
transform 1 0 9844 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_107
timestamp 0
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 0
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_138
timestamp 0
transform 1 0 13800 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_150
timestamp 0
transform 1 0 14904 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_173
timestamp 0
transform 1 0 17020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_185
timestamp 0
transform 1 0 18124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_197
timestamp 0
transform 1 0 19228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_209
timestamp 0
transform 1 0 20332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_221
timestamp 0
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_37
timestamp 0
transform 1 0 4508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_41
timestamp 0
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_48
timestamp 0
transform 1 0 5520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_57
timestamp 0
transform 1 0 6348 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_62
timestamp 0
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_72
timestamp 0
transform 1 0 7728 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_79
timestamp 0
transform 1 0 8372 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 0
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_85
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_90
timestamp 0
transform 1 0 9384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_97
timestamp 0
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_104
timestamp 0
transform 1 0 10672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_111
timestamp 0
transform 1 0 11316 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_141
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_149
timestamp 0
transform 1 0 14812 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_153
timestamp 0
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_167
timestamp 0
transform 1 0 16468 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_184
timestamp 0
transform 1 0 18032 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_191
timestamp 0
transform 1 0 18676 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 0
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_202
timestamp 0
transform 1 0 19688 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_214
timestamp 0
transform 1 0 20792 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_222
timestamp 0
transform 1 0 21528 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_225
timestamp 0
transform 1 0 21804 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 5520 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform 1 0 8464 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform -1 0 9384 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 11040 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform -1 0 15640 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 0
transform -1 0 13984 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 0
transform 1 0 18768 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 0
transform 1 0 21804 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 0
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 0
transform 1 0 21804 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 0
transform -1 0 22080 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform -1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 0
transform -1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 0
transform 1 0 21804 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 0
transform 1 0 21804 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 0
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 0
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 0
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 0
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 0
transform -1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 0
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 0
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 0
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 0
transform 1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 0
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 0
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 0
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 0
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 0
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 0
transform 1 0 4600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 0
transform -1 0 6808 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 0
transform -1 0 10028 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 0
transform 1 0 10396 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 0
transform -1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 0
transform -1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 0
transform 1 0 17756 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 0
transform -1 0 19688 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 0
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 0
transform 1 0 21804 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 0
transform 1 0 21804 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 0
transform -1 0 22080 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 0
transform -1 0 22080 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 0
transform -1 0 22080 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 0
transform 1 0 21804 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 0
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 0
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 0
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 0
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 0
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 0
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 0
transform -1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 0
transform -1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 0
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 0
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 0
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input66
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 0
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 0
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 0
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 0
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 0
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 0
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 0
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 0
transform 1 0 7176 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 0
transform 1 0 7820 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 0
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 0
transform 1 0 18124 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 0
transform -1 0 12604 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 0
transform 1 0 14260 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 0
transform 1 0 16652 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 0
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 0
transform 1 0 17204 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 0
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 0
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 0
transform -1 0 12052 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 0
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 0
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 0
transform 1 0 21712 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 0
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 0
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 0
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 0
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 0
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 0
transform 1 0 21712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 0
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 0
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 0
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 0
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 0
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 0
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output104
timestamp 0
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 22356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 22356 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 22356 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 22356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 22356 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 22356 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 22356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 22356 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 22356 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 22356 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 22356 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 22356 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 22356 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 22356 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 22356 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 22356 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 22356 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 22356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 22356 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 22356 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 22356 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 22356 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 22356 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 22356 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 0
transform -1 0 22356 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 0
transform -1 0 22356 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 0
transform -1 0 22356 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 0
transform -1 0 22356 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 0
transform -1 0 22356 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 0
transform -1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 0
transform -1 0 22356 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 0
transform -1 0 22356 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp 0
transform -1 0 17020 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer4
timestamp 0
transform 1 0 14444 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer5
timestamp 0
transform -1 0 14720 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer6
timestamp 0
transform -1 0 17940 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer7
timestamp 0
transform -1 0 15364 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer8
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9
timestamp 0
transform -1 0 20056 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer10
timestamp 0
transform 1 0 16928 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer11
timestamp 0
transform 1 0 18492 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_86
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_87
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_88
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_90
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_91
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_92
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_93
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_95
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_96
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_97
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_101
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_110
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_111
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_114
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_115
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_116
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_118
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_119
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_120
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_121
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_122
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_123
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_124
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_125
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_127
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_128
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_129
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_130
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_131
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_132
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_133
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_134
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_135
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_136
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_137
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_138
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_139
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_140
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_141
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_142
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_143
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_144
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_145
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_146
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_147
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_148
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_149
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_150
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_151
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_152
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_153
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_154
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_155
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_156
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_157
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_158
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_159
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_160
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_161
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_162
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_163
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_164
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_165
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_166
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_167
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_168
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_169
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_170
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_171
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_172
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_173
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_174
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_175
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_176
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_177
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_178
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_179
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_180
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_181
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_182
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_183
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_184
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_185
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_186
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_187
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_188
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_189
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_190
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_191
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_192
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_193
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_194
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_195
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_196
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_197
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_198
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_199
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_200
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_201
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_202
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_203
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_204
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_205
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_206
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_207
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_208
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_209
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_210
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_211
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_212
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_213
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_214
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_215
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_216
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_217
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_218
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_219
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_220
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_221
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_222
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_223
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_224
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_225
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_226
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_227
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_228
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_229
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_230
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_231
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_232
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_233
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_234
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_235
timestamp 0
transform 1 0 6256 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_236
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_237
timestamp 0
transform 1 0 11408 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_238
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_239
timestamp 0
transform 1 0 16560 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 0
transform 1 0 21712 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire105
timestamp 0
transform -1 0 7728 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire106
timestamp 0
transform -1 0 8924 0 -1 16320
box -38 -48 314 592
<< labels >>
rlabel metal1 s 11730 22848 11730 22848 4 VGND
rlabel metal1 s 11730 23392 11730 23392 4 VPWR
rlabel metal1 s 13754 6222 13754 6222 4 _0030_
rlabel metal1 s 15548 16422 15548 16422 4 _0032_
rlabel metal2 s 12742 9860 12742 9860 4 _0033_
rlabel metal2 s 12466 8942 12466 8942 4 _0034_
rlabel metal1 s 8142 17510 8142 17510 4 _0035_
rlabel metal1 s 12466 10132 12466 10132 4 _0036_
rlabel metal1 s 13478 18122 13478 18122 4 _0037_
rlabel metal1 s 13800 9894 13800 9894 4 _0038_
rlabel metal2 s 12834 9826 12834 9826 4 _0039_
rlabel metal2 s 7498 15436 7498 15436 4 _0040_
rlabel metal1 s 12834 9928 12834 9928 4 _0041_
rlabel metal1 s 8418 8942 8418 8942 4 _0043_
rlabel metal1 s 6210 15878 6210 15878 4 _0044_
rlabel metal1 s 6647 17510 6647 17510 4 _0045_
rlabel metal2 s 6210 17612 6210 17612 4 _0046_
rlabel metal2 s 7406 18700 7406 18700 4 _0047_
rlabel metal2 s 7590 18428 7590 18428 4 _0048_
rlabel metal2 s 6762 16320 6762 16320 4 _0049_
rlabel metal1 s 15640 17170 15640 17170 4 _0050_
rlabel metal1 s 13754 19380 13754 19380 4 _0051_
rlabel metal1 s 14076 19346 14076 19346 4 _0052_
rlabel metal2 s 15870 18870 15870 18870 4 _0053_
rlabel metal2 s 8418 7276 8418 7276 4 _0054_
rlabel metal1 s 16146 18190 16146 18190 4 _0055_
rlabel metal1 s 15962 16694 15962 16694 4 _0056_
rlabel metal2 s 15410 16354 15410 16354 4 _0057_
rlabel metal1 s 13340 15130 13340 15130 4 _0058_
rlabel metal1 s 15180 9078 15180 9078 4 _0059_
rlabel metal1 s 17204 10030 17204 10030 4 _0060_
rlabel metal2 s 16882 9758 16882 9758 4 _0061_
rlabel metal1 s 16054 7854 16054 7854 4 _0062_
rlabel metal1 s 16928 8466 16928 8466 4 _0063_
rlabel metal1 s 15180 7378 15180 7378 4 _0064_
rlabel metal2 s 7682 6902 7682 6902 4 _0065_
rlabel metal1 s 14306 7378 14306 7378 4 _0066_
rlabel metal1 s 15962 8908 15962 8908 4 _0067_
rlabel metal1 s 6762 7854 6762 7854 4 _0068_
rlabel metal2 s 7222 7684 7222 7684 4 _0069_
rlabel metal1 s 5658 10064 5658 10064 4 _0070_
rlabel metal1 s 6716 9554 6716 9554 4 _0071_
rlabel metal2 s 8234 9452 8234 9452 4 _0072_
rlabel metal1 s 7544 17578 7544 17578 4 _0073_
rlabel metal2 s 6486 15028 6486 15028 4 _0074_
rlabel metal1 s 11270 8908 11270 8908 4 _0079_
rlabel metal2 s 10442 8330 10442 8330 4 _0080_
rlabel metal1 s 8832 8602 8832 8602 4 _0081_
rlabel metal1 s 10541 8466 10541 8466 4 _0082_
rlabel metal1 s 10350 7922 10350 7922 4 _0084_
rlabel metal1 s 9246 8058 9246 8058 4 _0085_
rlabel metal2 s 9982 7582 9982 7582 4 _0086_
rlabel metal2 s 10166 7582 10166 7582 4 _0087_
rlabel metal1 s 10396 5746 10396 5746 4 _0088_
rlabel metal2 s 11270 8160 11270 8160 4 _0090_
rlabel metal1 s 12006 8058 12006 8058 4 _0094_
rlabel metal2 s 11546 8772 11546 8772 4 _0105_
rlabel metal2 s 12650 7650 12650 7650 4 _0108_
rlabel metal1 s 9568 8602 9568 8602 4 _0111_
rlabel metal1 s 12581 5542 12581 5542 4 _0120_
rlabel metal1 s 11914 5338 11914 5338 4 _0121_
rlabel metal1 s 13110 7514 13110 7514 4 _0122_
rlabel metal1 s 12788 7378 12788 7378 4 _0123_
rlabel metal1 s 12627 7310 12627 7310 4 _0125_
rlabel metal1 s 12926 7446 12926 7446 4 _0126_
rlabel metal2 s 13018 5882 13018 5882 4 _0127_
rlabel metal2 s 13202 5882 13202 5882 4 _0128_
rlabel metal1 s 13064 6290 13064 6290 4 _0131_
rlabel metal2 s 12742 8738 12742 8738 4 _0146_
rlabel metal1 s 12604 8058 12604 8058 4 _0152_
rlabel metal1 s 3105 15402 3105 15402 4 _0161_
rlabel metal1 s 2047 15130 2047 15130 4 _0162_
rlabel metal1 s 4094 15130 4094 15130 4 _0163_
rlabel metal1 s 3082 14960 3082 14960 4 _0164_
rlabel metal1 s 3174 15028 3174 15028 4 _0166_
rlabel metal2 s 4094 15708 4094 15708 4 _0167_
rlabel metal1 s 3174 15130 3174 15130 4 _0168_
rlabel metal1 s 4232 16082 4232 16082 4 _0169_
rlabel metal1 s 4048 17646 4048 17646 4 _0170_
rlabel metal1 s 4232 14994 4232 14994 4 _0172_
rlabel metal2 s 5658 15504 5658 15504 4 _0176_
rlabel metal1 s 4876 14926 4876 14926 4 _0178_
rlabel metal2 s 5474 15708 5474 15708 4 _0187_
rlabel metal1 s 5060 15402 5060 15402 4 _0193_
rlabel metal1 s 2507 17850 2507 17850 4 _0202_
rlabel metal2 s 1978 17884 1978 17884 4 _0203_
rlabel metal2 s 3358 18496 3358 18496 4 _0204_
rlabel metal1 s 3772 18734 3772 18734 4 _0205_
rlabel metal1 s 3588 18802 3588 18802 4 _0207_
rlabel metal1 s 3036 18394 3036 18394 4 _0208_
rlabel metal1 s 4002 18666 4002 18666 4 _0209_
rlabel metal1 s 4600 18326 4600 18326 4 _0210_
rlabel metal1 s 5106 19346 5106 19346 4 _0211_
rlabel metal1 s 3772 17714 3772 17714 4 _0213_
rlabel metal1 s 4830 17578 4830 17578 4 _0217_
rlabel metal1 s 5750 17510 5750 17510 4 _0228_
rlabel metal2 s 6026 17884 6026 17884 4 _0234_
rlabel metal1 s 5497 21522 5497 21522 4 _0243_
rlabel metal2 s 4554 21148 4554 21148 4 _0244_
rlabel metal1 s 6026 19924 6026 19924 4 _0245_
rlabel metal1 s 5612 20842 5612 20842 4 _0246_
rlabel metal2 s 5658 20179 5658 20179 4 _0248_
rlabel metal1 s 5382 20570 5382 20570 4 _0249_
rlabel metal1 s 5060 20502 5060 20502 4 _0250_
rlabel metal1 s 5658 20026 5658 20026 4 _0251_
rlabel metal1 s 7406 20434 7406 20434 4 _0252_
rlabel metal1 s 5106 19856 5106 19856 4 _0254_
rlabel metal2 s 5934 18938 5934 18938 4 _0258_
rlabel metal2 s 5658 18496 5658 18496 4 _0269_
rlabel metal2 s 5750 19312 5750 19312 4 _0275_
rlabel metal1 s 8188 21658 8188 21658 4 _0284_
rlabel metal1 s 8211 22678 8211 22678 4 _0285_
rlabel metal1 s 8004 21930 8004 21930 4 _0286_
rlabel metal1 s 8556 21522 8556 21522 4 _0287_
rlabel metal2 s 8602 21726 8602 21726 4 _0289_
rlabel metal1 s 7590 21998 7590 21998 4 _0290_
rlabel metal2 s 8326 21114 8326 21114 4 _0291_
rlabel metal1 s 7912 20842 7912 20842 4 _0292_
rlabel metal2 s 9338 20604 9338 20604 4 _0293_
rlabel metal1 s 7268 20978 7268 20978 4 _0295_
rlabel metal2 s 7590 20026 7590 20026 4 _0299_
rlabel metal2 s 7314 19584 7314 19584 4 _0310_
rlabel metal2 s 7406 20672 7406 20672 4 _0316_
rlabel metal1 s 11385 19482 11385 19482 4 _0325_
rlabel metal1 s 11247 20434 11247 20434 4 _0326_
rlabel metal1 s 10120 18938 10120 18938 4 _0327_
rlabel metal1 s 10764 19958 10764 19958 4 _0328_
rlabel metal2 s 10442 19992 10442 19992 4 _0330_
rlabel metal1 s 10672 19482 10672 19482 4 _0331_
rlabel metal1 s 9982 19414 9982 19414 4 _0332_
rlabel metal1 s 10350 20366 10350 20366 4 _0333_
rlabel metal1 s 10764 17714 10764 17714 4 _0334_
rlabel metal1 s 9568 19890 9568 19890 4 _0336_
rlabel metal2 s 8786 19686 8786 19686 4 _0340_
rlabel metal2 s 8418 18972 8418 18972 4 _0351_
rlabel metal1 s 9062 18734 9062 18734 4 _0357_
rlabel metal1 s 11339 16082 11339 16082 4 _0366_
rlabel metal1 s 10764 15538 10764 15538 4 _0367_
rlabel metal1 s 10120 16422 10120 16422 4 _0368_
rlabel metal2 s 10534 16864 10534 16864 4 _0369_
rlabel metal1 s 10764 17034 10764 17034 4 _0371_
rlabel metal1 s 9982 16660 9982 16660 4 _0372_
rlabel metal1 s 11132 17306 11132 17306 4 _0373_
rlabel metal1 s 11224 17646 11224 17646 4 _0374_
rlabel metal1 s 12558 17646 12558 17646 4 _0375_
rlabel metal2 s 10166 17408 10166 17408 4 _0377_
rlabel metal2 s 8878 17510 8878 17510 4 _0381_
rlabel metal2 s 8326 16796 8326 16796 4 _0392_
rlabel metal1 s 8878 16422 8878 16422 4 _0398_
rlabel metal1 s 13501 16218 13501 16218 4 _0407_
rlabel metal1 s 12811 16218 12811 16218 4 _0408_
rlabel metal1 s 13708 17170 13708 17170 4 _0409_
rlabel metal2 s 12926 17952 12926 17952 4 _0410_
rlabel metal1 s 12788 17646 12788 17646 4 _0412_
rlabel metal1 s 13432 17238 13432 17238 4 _0413_
rlabel metal1 s 13156 18258 13156 18258 4 _0414_
rlabel metal1 s 12834 17850 12834 17850 4 _0415_
rlabel metal1 s 13340 19346 13340 19346 4 _0416_
rlabel metal1 s 12834 17782 12834 17782 4 _0418_
rlabel metal1 s 15410 17680 15410 17680 4 _0422_
rlabel metal1 s 15226 17306 15226 17306 4 _0433_
rlabel metal1 s 14766 17238 14766 17238 4 _0439_
rlabel metal2 s 14145 22066 14145 22066 4 _0448_
rlabel metal1 s 13363 22746 13363 22746 4 _0449_
rlabel metal1 s 13524 21930 13524 21930 4 _0450_
rlabel metal1 s 12604 21454 12604 21454 4 _0451_
rlabel metal1 s 12742 21522 12742 21522 4 _0453_
rlabel metal1 s 12742 21998 12742 21998 4 _0454_
rlabel metal2 s 13478 21114 13478 21114 4 _0455_
rlabel metal2 s 13662 20672 13662 20672 4 _0456_
rlabel metal1 s 14628 20910 14628 20910 4 _0457_
rlabel metal2 s 13202 19856 13202 19856 4 _0459_
rlabel metal1 s 13386 19278 13386 19278 4 _0463_
rlabel metal1 s 12650 19754 12650 19754 4 _0474_
rlabel metal1 s 12604 19822 12604 19822 4 _0480_
rlabel metal1 s 15755 22746 15755 22746 4 _0489_
rlabel metal1 s 16169 22610 16169 22610 4 _0490_
rlabel metal1 s 14996 21930 14996 21930 4 _0491_
rlabel metal2 s 16146 21794 16146 21794 4 _0492_
rlabel metal1 s 15226 22066 15226 22066 4 _0494_
rlabel metal2 s 15962 21760 15962 21760 4 _0495_
rlabel metal1 s 15916 20842 15916 20842 4 _0496_
rlabel metal1 s 15870 20910 15870 20910 4 _0497_
rlabel metal2 s 17158 20672 17158 20672 4 _0498_
rlabel metal1 s 15456 21046 15456 21046 4 _0500_
rlabel metal2 s 15226 20026 15226 20026 4 _0504_
rlabel metal2 s 14766 19584 14766 19584 4 _0515_
rlabel metal2 s 14674 20672 14674 20672 4 _0521_
rlabel metal1 s 19941 20434 19941 20434 4 _0530_
rlabel metal1 s 19941 20774 19941 20774 4 _0531_
rlabel metal1 s 18308 20570 18308 20570 4 _0532_
rlabel metal1 s 18400 20910 18400 20910 4 _0533_
rlabel metal1 s 18722 20298 18722 20298 4 _0535_
rlabel metal1 s 18584 20570 18584 20570 4 _0536_
rlabel metal2 s 18906 20026 18906 20026 4 _0537_
rlabel metal1 s 18676 19822 18676 19822 4 _0538_
rlabel metal1 s 18492 17646 18492 17646 4 _0539_
rlabel metal1 s 17572 20366 17572 20366 4 _0541_
rlabel metal2 s 16790 20026 16790 20026 4 _0545_
rlabel metal2 s 17158 19584 17158 19584 4 _0556_
rlabel metal2 s 17066 19856 17066 19856 4 _0562_
rlabel metal1 s 11753 3706 11753 3706 4 _0571_
rlabel metal1 s 9913 3162 9913 3162 4 _0572_
rlabel metal2 s 10166 4386 10166 4386 4 _0573_
rlabel metal2 s 10810 4318 10810 4318 4 _0574_
rlabel metal1 s 9568 4114 9568 4114 4 _0576_
rlabel metal1 s 10028 4250 10028 4250 4 _0577_
rlabel metal1 s 9338 4794 9338 4794 4 _0578_
rlabel metal1 s 10258 5270 10258 5270 4 _0579_
rlabel metal1 s 9108 5134 9108 5134 4 _0580_
rlabel metal2 s 10074 5270 10074 5270 4 _0582_
rlabel metal2 s 9798 6086 9798 6086 4 _0586_
rlabel metal1 s 9522 6426 9522 6426 4 _0597_
rlabel metal2 s 9522 5508 9522 5508 4 _0603_
rlabel metal1 s 20861 17510 20861 17510 4 _0612_
rlabel metal1 s 20677 18258 20677 18258 4 _0613_
rlabel metal2 s 19366 17816 19366 17816 4 _0614_
rlabel metal1 s 19320 17170 19320 17170 4 _0615_
rlabel metal1 s 19918 18360 19918 18360 4 _0617_
rlabel metal1 s 19366 18258 19366 18258 4 _0618_
rlabel metal1 s 18998 17306 18998 17306 4 _0619_
rlabel metal2 s 18814 17442 18814 17442 4 _0620_
rlabel metal2 s 18722 17035 18722 17035 4 _0621_
rlabel metal1 s 18814 17714 18814 17714 4 _0623_
rlabel metal2 s 18078 18054 18078 18054 4 _0627_
rlabel metal1 s 17526 18394 17526 18394 4 _0638_
rlabel metal1 s 17986 18326 17986 18326 4 _0644_
rlabel metal2 s 21206 15232 21206 15232 4 _0653_
rlabel metal2 s 20401 14586 20401 14586 4 _0654_
rlabel metal2 s 19274 14790 19274 14790 4 _0655_
rlabel metal1 s 19642 14892 19642 14892 4 _0656_
rlabel metal1 s 19550 15028 19550 15028 4 _0658_
rlabel metal1 s 18032 15062 18032 15062 4 _0659_
rlabel metal1 s 18768 14042 18768 14042 4 _0660_
rlabel metal1 s 19044 14382 19044 14382 4 _0661_
rlabel metal1 s 17158 14382 17158 14382 4 _0662_
rlabel metal1 s 19366 15504 19366 15504 4 _0664_
rlabel metal2 s 18446 15878 18446 15878 4 _0668_
rlabel metal1 s 17894 16218 17894 16218 4 _0679_
rlabel metal2 s 18354 15606 18354 15606 4 _0685_
rlabel metal1 s 17365 13906 17365 13906 4 _0694_
rlabel metal1 s 15985 13158 15985 13158 4 _0695_
rlabel metal1 s 16100 14382 16100 14382 4 _0696_
rlabel metal1 s 17480 14314 17480 14314 4 _0697_
rlabel metal1 s 17434 14380 17434 14380 4 _0699_
rlabel metal1 s 16560 14314 16560 14314 4 _0700_
rlabel metal1 s 15870 13906 15870 13906 4 _0701_
rlabel metal1 s 16008 13974 16008 13974 4 _0702_
rlabel metal2 s 14674 14212 14674 14212 4 _0703_
rlabel metal2 s 15502 14756 15502 14756 4 _0705_
rlabel metal1 s 16238 14926 16238 14926 4 _0709_
rlabel metal2 s 15778 15844 15778 15844 4 _0720_
rlabel metal1 s 15640 14586 15640 14586 4 _0726_
rlabel metal2 s 12581 12410 12581 12410 4 _0735_
rlabel metal2 s 12121 12954 12121 12954 4 _0736_
rlabel metal1 s 12006 13498 12006 13498 4 _0737_
rlabel metal2 s 11546 13668 11546 13668 4 _0738_
rlabel metal2 s 12834 13022 12834 13022 4 _0740_
rlabel metal1 s 12374 13906 12374 13906 4 _0741_
rlabel metal1 s 13570 12818 13570 12818 4 _0742_
rlabel metal1 s 13616 12886 13616 12886 4 _0743_
rlabel metal1 s 14674 12614 14674 12614 4 _0744_
rlabel metal1 s 13754 13294 13754 13294 4 _0746_
rlabel metal2 s 13386 14042 13386 14042 4 _0750_
rlabel metal2 s 13110 14756 13110 14756 4 _0761_
rlabel metal2 s 13018 14518 13018 14518 4 _0767_
rlabel metal1 s 15617 11050 15617 11050 4 _0776_
rlabel metal1 s 14030 11118 14030 11118 4 _0777_
rlabel metal2 s 14674 10234 14674 10234 4 _0778_
rlabel metal1 s 15088 10982 15088 10982 4 _0779_
rlabel metal1 s 14674 10982 14674 10982 4 _0781_
rlabel metal1 s 14950 10098 14950 10098 4 _0782_
rlabel metal1 s 14904 11322 14904 11322 4 _0783_
rlabel metal1 s 15916 11798 15916 11798 4 _0784_
rlabel metal1 s 16606 11186 16606 11186 4 _0785_
rlabel metal1 s 14628 11526 14628 11526 4 _0787_
rlabel metal2 s 15502 9724 15502 9724 4 _0791_
rlabel metal1 s 14858 8874 14858 8874 4 _0802_
rlabel metal2 s 14674 9418 14674 9418 4 _0808_
rlabel metal1 s 20217 12410 20217 12410 4 _0817_
rlabel metal1 s 19596 12750 19596 12750 4 _0818_
rlabel metal1 s 18492 12206 18492 12206 4 _0819_
rlabel metal1 s 19044 12750 19044 12750 4 _0820_
rlabel metal1 s 19090 12682 19090 12682 4 _0822_
rlabel metal2 s 18354 11968 18354 11968 4 _0823_
rlabel metal2 s 18492 11050 18492 11050 4 _0824_
rlabel metal1 s 18768 11118 18768 11118 4 _0825_
rlabel metal1 s 18814 10098 18814 10098 4 _0826_
rlabel metal2 s 17710 11730 17710 11730 4 _0828_
rlabel metal2 s 18170 11526 18170 11526 4 _0832_
rlabel metal1 s 17342 11866 17342 11866 4 _0843_
rlabel metal1 s 17572 11798 17572 11798 4 _0849_
rlabel metal1 s 21137 9690 21137 9690 4 _0858_
rlabel metal2 s 20562 10268 20562 10268 4 _0859_
rlabel metal1 s 20148 9690 20148 9690 4 _0860_
rlabel metal1 s 19688 10642 19688 10642 4 _0861_
rlabel metal1 s 19504 10574 19504 10574 4 _0863_
rlabel metal1 s 19596 10098 19596 10098 4 _0864_
rlabel metal2 s 20194 9605 20194 9605 4 _0865_
rlabel metal1 s 19366 9146 19366 9146 4 _0866_
rlabel metal2 s 20010 8908 20010 8908 4 _0867_
rlabel metal2 s 18814 9248 18814 9248 4 _0869_
rlabel metal1 s 18308 9486 18308 9486 4 _0873_
rlabel metal1 s 17526 9894 17526 9894 4 _0884_
rlabel metal1 s 18262 9962 18262 9962 4 _0890_
rlabel metal2 s 20930 7004 20930 7004 4 _0899_
rlabel metal1 s 20953 7378 20953 7378 4 _0900_
rlabel metal1 s 19228 7514 19228 7514 4 _0901_
rlabel metal1 s 19550 7276 19550 7276 4 _0902_
rlabel metal1 s 19412 7378 19412 7378 4 _0904_
rlabel metal2 s 19918 7344 19918 7344 4 _0905_
rlabel metal1 s 19642 6426 19642 6426 4 _0906_
rlabel metal1 s 18768 7446 18768 7446 4 _0907_
rlabel metal1 s 18814 6834 18814 6834 4 _0908_
rlabel metal1 s 19136 7922 19136 7922 4 _0910_
rlabel metal1 s 17848 7786 17848 7786 4 _0914_
rlabel metal1 s 17066 7718 17066 7718 4 _0925_
rlabel metal1 s 17158 7786 17158 7786 4 _0931_
rlabel metal1 s 20677 4454 20677 4454 4 _0940_
rlabel metal2 s 19297 3706 19297 3706 4 _0941_
rlabel metal2 s 17710 4998 17710 4998 4 _0942_
rlabel metal1 s 19458 4488 19458 4488 4 _0943_
rlabel metal1 s 19412 4590 19412 4590 4 _0945_
rlabel metal2 s 19274 4930 19274 4930 4 _0946_
rlabel metal1 s 18584 4522 18584 4522 4 _0947_
rlabel metal1 s 18768 4590 18768 4590 4 _0948_
rlabel metal2 s 17894 4964 17894 4964 4 _0949_
rlabel metal2 s 18906 5406 18906 5406 4 _0951_
rlabel metal2 s 18446 6426 18446 6426 4 _0955_
rlabel metal1 s 17526 6630 17526 6630 4 _0966_
rlabel metal2 s 18262 6018 18262 6018 4 _0972_
rlabel metal1 s 17940 3162 17940 3162 4 _0981_
rlabel metal1 s 16813 2958 16813 2958 4 _0982_
rlabel metal2 s 17066 3910 17066 3910 4 _0983_
rlabel metal2 s 16882 3332 16882 3332 4 _0984_
rlabel metal1 s 16606 3570 16606 3570 4 _0986_
rlabel metal1 s 16330 3978 16330 3978 4 _0987_
rlabel metal1 s 16790 3706 16790 3706 4 _0988_
rlabel metal1 s 17158 4488 17158 4488 4 _0989_
rlabel metal1 s 14950 4658 14950 4658 4 _0990_
rlabel metal2 s 16698 4318 16698 4318 4 _0992_
rlabel metal1 s 17158 5134 17158 5134 4 _0996_
rlabel metal2 s 16698 6528 16698 6528 4 _1007_
rlabel metal1 s 16652 3910 16652 3910 4 _1013_
rlabel metal1 s 7797 3026 7797 3026 4 _1022_
rlabel metal1 s 7084 2482 7084 2482 4 _1023_
rlabel metal2 s 7498 4352 7498 4352 4 _1024_
rlabel metal1 s 6854 4046 6854 4046 4 _1025_
rlabel metal1 s 6854 3434 6854 3434 4 _1027_
rlabel metal2 s 7406 3876 7406 3876 4 _1028_
rlabel metal1 s 6348 3706 6348 3706 4 _1029_
rlabel metal1 s 7728 5270 7728 5270 4 _1030_
rlabel metal1 s 6394 5134 6394 5134 4 _1031_
rlabel metal1 s 7406 5134 7406 5134 4 _1033_
rlabel metal2 s 7958 5338 7958 5338 4 _1037_
rlabel metal2 s 7590 6052 7590 6052 4 _1048_
rlabel metal1 s 7774 3978 7774 3978 4 _1054_
rlabel metal1 s 14421 2890 14421 2890 4 _1063_
rlabel metal2 s 14306 3264 14306 3264 4 _1064_
rlabel metal1 s 13662 3706 13662 3706 4 _1065_
rlabel metal1 s 14214 3434 14214 3434 4 _1066_
rlabel metal2 s 13570 3298 13570 3298 4 _1068_
rlabel metal1 s 13984 3706 13984 3706 4 _1069_
rlabel metal1 s 13432 4250 13432 4250 4 _1070_
rlabel metal2 s 13754 4862 13754 4862 4 _1071_
rlabel metal1 s 14260 5202 14260 5202 4 _1074_
rlabel metal1 s 14950 4794 14950 4794 4 _1078_
rlabel metal1 s 14582 5882 14582 5882 4 _1089_
rlabel metal1 s 14674 3978 14674 3978 4 _1095_
rlabel metal1 s 5313 3978 5313 3978 4 _1104_
rlabel metal2 s 4094 5882 4094 5882 4 _1105_
rlabel metal1 s 4232 5338 4232 5338 4 _1106_
rlabel metal1 s 4048 5134 4048 5134 4 _1107_
rlabel metal1 s 4094 5814 4094 5814 4 _1109_
rlabel metal1 s 4784 5338 4784 5338 4 _1110_
rlabel metal1 s 3634 5882 3634 5882 4 _1111_
rlabel metal1 s 4646 6358 4646 6358 4 _1112_
rlabel metal1 s 4922 7310 4922 7310 4 _1113_
rlabel metal1 s 5428 5746 5428 5746 4 _1115_
rlabel metal2 s 6118 6086 6118 6086 4 _1119_
rlabel metal1 s 6256 6426 6256 6426 4 _1130_
rlabel metal2 s 5290 6562 5290 6562 4 _1136_
rlabel metal2 s 2622 7616 2622 7616 4 _1145_
rlabel metal1 s 1955 7514 1955 7514 4 _1146_
rlabel metal1 s 4232 7854 4232 7854 4 _1147_
rlabel metal1 s 3220 8466 3220 8466 4 _1148_
rlabel metal1 s 3220 7922 3220 7922 4 _1150_
rlabel metal1 s 4232 7922 4232 7922 4 _1151_
rlabel metal1 s 3818 8058 3818 8058 4 _1152_
rlabel metal1 s 4232 8466 4232 8466 4 _1153_
rlabel metal1 s 4232 9486 4232 9486 4 _1154_
rlabel metal1 s 4278 7378 4278 7378 4 _1156_
rlabel metal2 s 5566 8092 5566 8092 4 _1160_
rlabel metal2 s 5382 7616 5382 7616 4 _1171_
rlabel metal1 s 5290 7446 5290 7446 4 _1177_
rlabel metal2 s 2346 10404 2346 10404 4 _1186_
rlabel metal2 s 2254 10812 2254 10812 4 _1187_
rlabel metal1 s 2185 10778 2185 10778 4 _1188_
rlabel metal1 s 2162 10574 2162 10574 4 _1189_
rlabel metal1 s 2714 10132 2714 10132 4 _1191_
rlabel metal1 s 3220 10778 3220 10778 4 _1192_
rlabel metal1 s 3726 10234 3726 10234 4 _1193_
rlabel metal1 s 4784 9622 4784 9622 4 _1194_
rlabel metal1 s 6854 10642 6854 10642 4 _1195_
rlabel metal1 s 4232 10098 4232 10098 4 _1197_
rlabel metal2 s 4554 10438 4554 10438 4 _1201_
rlabel metal2 s 4922 10268 4922 10268 4 _1212_
rlabel metal2 s 5014 10268 5014 10268 4 _1218_
rlabel metal1 s 7705 12070 7705 12070 4 _1227_
rlabel metal1 s 7613 12818 7613 12818 4 _1228_
rlabel metal1 s 7038 11866 7038 11866 4 _1229_
rlabel metal2 s 7038 11628 7038 11628 4 _1230_
rlabel metal1 s 6762 12342 6762 12342 4 _1232_
rlabel metal1 s 7820 11798 7820 11798 4 _1233_
rlabel metal2 s 7682 11322 7682 11322 4 _1234_
rlabel metal1 s 7912 10710 7912 10710 4 _1235_
rlabel metal2 s 8602 11458 8602 11458 4 _1236_
rlabel metal1 s 7268 10642 7268 10642 4 _1238_
rlabel metal1 s 7268 8942 7268 8942 4 _1242_
rlabel metal1 s 6578 8874 6578 8874 4 _1253_
rlabel metal2 s 6394 10234 6394 10234 4 _1259_
rlabel metal2 s 11661 10778 11661 10778 4 _1268_
rlabel metal2 s 12075 10778 12075 10778 4 _1269_
rlabel metal2 s 10626 11322 10626 11322 4 _1270_
rlabel metal1 s 11086 11254 11086 11254 4 _1271_
rlabel metal1 s 10350 11730 10350 11730 4 _1273_
rlabel metal1 s 10764 10234 10764 10234 4 _1274_
rlabel metal1 s 9890 12138 9890 12138 4 _1275_
rlabel metal2 s 8970 12002 8970 12002 4 _1276_
rlabel metal2 s 8694 14076 8694 14076 4 _1277_
rlabel metal1 s 8970 11662 8970 11662 4 _1279_
rlabel metal2 s 9430 11322 9430 11322 4 _1283_
rlabel metal1 s 9154 10778 9154 10778 4 _1294_
rlabel metal1 s 9706 10710 9706 10710 4 _1300_
rlabel metal1 s 10557 13906 10557 13906 4 _1309_
rlabel metal2 s 10350 13532 10350 13532 4 _1310_
rlabel metal2 s 9430 14790 9430 14790 4 _1311_
rlabel metal1 s 9292 13838 9292 13838 4 _1312_
rlabel metal1 s 9430 13430 9430 13430 4 _1314_
rlabel metal1 s 8878 14586 8878 14586 4 _1315_
rlabel metal1 s 9384 13226 9384 13226 4 _1316_
rlabel metal1 s 9890 13294 9890 13294 4 _1317_
rlabel metal1 s 6394 13906 6394 13906 4 _1318_
rlabel metal1 s 9752 13838 9752 13838 4 _1320_
rlabel metal1 s 8234 13838 8234 13838 4 _1324_
rlabel metal2 s 7774 15266 7774 15266 4 _1335_
rlabel metal1 s 8556 14858 8556 14858 4 _1341_
rlabel metal1 s 4715 12410 4715 12410 4 _1350_
rlabel metal1 s 4048 12750 4048 12750 4 _1351_
rlabel metal1 s 5382 13226 5382 13226 4 _1352_
rlabel metal1 s 5750 13328 5750 13328 4 _1353_
rlabel metal1 s 4278 13260 4278 13260 4 _1355_
rlabel metal1 s 5290 13294 5290 13294 4 _1356_
rlabel metal1 s 5060 12954 5060 12954 4 _1357_
rlabel metal1 s 5060 13974 5060 13974 4 _1358_
rlabel metal2 s 5934 13668 5934 13668 4 _1361_
rlabel metal2 s 6394 14042 6394 14042 4 _1365_
rlabel metal1 s 5934 14314 5934 14314 4 _1376_
rlabel metal1 s 5612 13498 5612 13498 4 _1382_
rlabel metal2 s 3266 1588 3266 1588 4 a[0]
rlabel metal3 s 1050 15028 1050 15028 4 a[10]
rlabel metal3 s 0 21768 800 21888 4 a[11]
port 5 nsew
rlabel metal2 s 5290 24021 5290 24021 4 a[12]
rlabel metal1 s 8556 23086 8556 23086 4 a[13]
rlabel metal1 s 9246 23086 9246 23086 4 a[14]
rlabel metal1 s 11040 23086 11040 23086 4 a[15]
rlabel metal2 s 15594 24021 15594 24021 4 a[16]
rlabel metal1 s 13662 23086 13662 23086 4 a[17]
rlabel metal2 s 18998 24021 18998 24021 4 a[18]
rlabel metal2 s 22034 20689 22034 20689 4 a[19]
rlabel metal2 s 10994 1588 10994 1588 4 a[1]
rlabel metal3 s 22034 19805 22034 19805 4 a[20]
rlabel metal2 s 22034 15895 22034 15895 4 a[21]
rlabel metal2 s 22034 19227 22034 19227 4 a[22]
rlabel metal2 s 22034 12563 22034 12563 4 a[23]
rlabel metal2 s 22034 11679 22034 11679 4 a[24]
rlabel metal3 s 22034 14365 22034 14365 4 a[25]
rlabel metal2 s 22034 5015 22034 5015 4 a[26]
rlabel metal2 s 22034 5593 22034 5593 4 a[27]
rlabel metal2 s 22034 4369 22034 4369 4 a[28]
rlabel metal2 s 20010 1588 20010 1588 4 a[29]
rlabel metal2 s 5198 1588 5198 1588 4 a[2]
rlabel metal2 s 17434 1588 17434 1588 4 a[30]
rlabel metal2 s 12282 1588 12282 1588 4 a[31]
rlabel metal2 s 4554 1027 4554 1027 4 a[3]
rlabel metal3 s 0 6128 800 6248 4 a[4]
port 29 nsew
rlabel metal3 s 0 7488 800 7608 4 a[5]
port 30 nsew
rlabel metal3 s 1188 10948 1188 10948 4 a[6]
rlabel metal2 s 11638 1588 11638 1588 4 a[7]
rlabel metal3 s 1050 13668 1050 13668 4 a[8]
rlabel metal3 s 1050 12308 1050 12308 4 a[9]
rlabel metal3 s 0 3408 800 3528 4 ainv
port 35 nsew
rlabel metal2 s 10350 1588 10350 1588 4 b[0]
rlabel metal3 s 0 16328 800 16448 4 b[10]
port 37 nsew
rlabel metal3 s 0 18368 800 18488 4 b[11]
port 38 nsew
rlabel metal2 s 4830 24021 4830 24021 4 b[12]
rlabel metal2 s 6578 24021 6578 24021 4 b[13]
rlabel metal1 s 9752 23086 9752 23086 4 b[14]
rlabel metal2 s 10442 24021 10442 24021 4 b[15]
rlabel metal2 s 15134 24021 15134 24021 4 b[16]
rlabel metal1 s 13202 23086 13202 23086 4 b[17]
rlabel metal1 s 17710 23086 17710 23086 4 b[18]
rlabel metal2 s 19458 24021 19458 24021 4 b[19]
rlabel metal2 s 9706 823 9706 823 4 b[1]
rlabel metal2 s 22034 18581 22034 18581 4 b[20]
rlabel metal2 s 22034 15249 22034 15249 4 b[21]
rlabel metal2 s 22034 16473 22034 16473 4 b[22]
rlabel metal2 s 22034 13787 22034 13787 4 b[23]
rlabel metal2 s 22034 11033 22034 11033 4 b[24]
rlabel metal2 s 22034 13141 22034 13141 4 b[25]
rlabel metal2 s 22034 10455 22034 10455 4 b[26]
rlabel metal2 s 22034 7123 22034 7123 4 b[27]
rlabel metal2 s 19366 1588 19366 1588 4 b[28]
rlabel metal2 s 18078 1588 18078 1588 4 b[29]
rlabel metal2 s 6486 1588 6486 1588 4 b[2]
rlabel metal2 s 14858 1027 14858 1027 4 b[30]
rlabel metal2 s 13570 1588 13570 1588 4 b[31]
rlabel metal3 s 0 4768 800 4888 4 b[3]
port 61 nsew
rlabel metal3 s 1188 6868 1188 6868 4 b[4]
rlabel metal3 s 1096 10268 1096 10268 4 b[5]
rlabel metal3 s 0 11568 800 11688 4 b[6]
port 64 nsew
rlabel metal2 s 3910 1588 3910 1588 4 b[7]
rlabel metal3 s 0 14288 800 14408 4 b[8]
port 66 nsew
rlabel metal3 s 0 12928 800 13048 4 b[9]
port 67 nsew
rlabel metal3 s 0 22448 800 22568 4 binv
port 68 nsew
rlabel metal2 s 9062 1588 9062 1588 4 cin
rlabel metal2 s 14214 1520 14214 1520 4 cout
rlabel metal1 s 3542 2516 3542 2516 4 net1
rlabel metal1 s 16376 23086 16376 23086 4 net10
rlabel metal1 s 2231 8942 2231 8942 4 net100
rlabel metal1 s 6762 2312 6762 2312 4 net101
rlabel metal1 s 7544 16422 7544 16422 4 net102
rlabel metal1 s 6210 15674 6210 15674 4 net103
rlabel metal1 s 13064 2414 13064 2414 4 net104
rlabel metal1 s 10304 14790 10304 14790 4 net105
rlabel metal2 s 12282 12444 12282 12444 4 net106
rlabel metal1 s 12834 8976 12834 8976 4 net107
rlabel metal2 s 16146 6596 16146 6596 4 net108
rlabel metal1 s 5704 18190 5704 18190 4 net109
rlabel metal1 s 21050 20434 21050 20434 4 net11
rlabel metal1 s 17388 19278 17388 19278 4 net110
rlabel metal1 s 9062 8466 9062 8466 4 net111
rlabel metal1 s 10258 11186 10258 11186 4 net112
rlabel metal2 s 13294 8194 13294 8194 4 net113
rlabel metal1 s 18400 11662 18400 11662 4 net114
rlabel metal2 s 4922 17884 4922 17884 4 net115
rlabel metal1 s 6348 18802 6348 18802 4 net116
rlabel metal1 s 18630 15980 18630 15980 4 net117
rlabel metal1 s 18814 18190 18814 18190 4 net118
rlabel metal1 s 5152 13906 5152 13906 4 net119
rlabel metal1 s 11671 3502 11671 3502 4 net12
rlabel metal1 s 1840 7922 1840 7922 4 net120
rlabel metal2 s 12558 11356 12558 11356 4 net121
rlabel metal2 s 4738 19414 4738 19414 4 net122
rlabel metal1 s 20240 20978 20240 20978 4 net123
rlabel metal1 s 2645 7922 2645 7922 4 net124
rlabel metal1 s 12466 12716 12466 12716 4 net125
rlabel metal1 s 5704 21454 5704 21454 4 net126
rlabel metal1 s 20700 17714 20700 17714 4 net127
rlabel metal1 s 15686 19822 15686 19822 4 net128
rlabel metal1 s 16974 19754 16974 19754 4 net129
rlabel metal1 s 21510 17646 21510 17646 4 net13
rlabel metal1 s 10350 6290 10350 6290 4 net130
rlabel metal2 s 18170 18564 18170 18564 4 net131
rlabel metal1 s 18722 16082 18722 16082 4 net132
rlabel metal2 s 16238 15708 16238 15708 4 net133
rlabel metal2 s 13570 14620 13570 14620 4 net134
rlabel metal2 s 15594 9180 15594 9180 4 net135
rlabel metal1 s 17940 11866 17940 11866 4 net136
rlabel metal1 s 18216 9554 18216 9554 4 net137
rlabel metal1 s 17664 7922 17664 7922 4 net138
rlabel metal1 s 18354 6766 18354 6766 4 net139
rlabel metal2 s 21114 15504 21114 15504 4 net14
rlabel metal1 s 16836 6222 16836 6222 4 net140
rlabel metal1 s 8050 5780 8050 5780 4 net141
rlabel metal2 s 14950 5916 14950 5916 4 net142
rlabel metal2 s 6854 6596 6854 6596 4 net143
rlabel metal2 s 5658 8092 5658 8092 4 net144
rlabel metal1 s 5152 10778 5152 10778 4 net145
rlabel metal1 s 7130 8806 7130 8806 4 net146
rlabel metal1 s 9706 11118 9706 11118 4 net147
rlabel metal1 s 8418 15130 8418 15130 4 net148
rlabel metal1 s 6854 14382 6854 14382 4 net149
rlabel metal1 s 21758 19482 21758 19482 4 net15
rlabel metal2 s 13386 8704 13386 8704 4 net150
rlabel metal1 s 5704 16218 5704 16218 4 net151
rlabel metal1 s 5152 17714 5152 17714 4 net152
rlabel metal1 s 6394 18734 6394 18734 4 net153
rlabel metal1 s 7866 19822 7866 19822 4 net154
rlabel metal1 s 8602 19278 8602 19278 4 net155
rlabel metal2 s 8970 17476 8970 17476 4 net156
rlabel metal1 s 15686 17646 15686 17646 4 net157
rlabel metal1 s 13570 19822 13570 19822 4 net158
rlabel metal2 s 2162 9894 2162 9894 4 net159
rlabel metal1 s 21850 12750 21850 12750 4 net16
rlabel metal1 s 4462 12716 4462 12716 4 net160
rlabel metal2 s 16514 14790 16514 14790 4 net161
rlabel metal1 s 15226 4590 15226 4590 4 net162
rlabel metal2 s 13754 14076 13754 14076 4 net163
rlabel metal1 s 17158 5202 17158 5202 4 net164
rlabel metal1 s 14628 10642 14628 10642 4 net165
rlabel metal2 s 18814 6460 18814 6460 4 net166
rlabel metal1 s 19182 7854 19182 7854 4 net167
rlabel metal1 s 17618 11118 17618 11118 4 net168
rlabel metal2 s 18906 9724 18906 9724 4 net169
rlabel metal2 s 15944 11118 15944 11118 4 net17
rlabel metal1 s 20516 12886 20516 12886 4 net18
rlabel metal2 s 21298 7616 21298 7616 4 net19
rlabel metal1 s 3194 15470 3194 15470 4 net2
rlabel metal1 s 21344 6630 21344 6630 4 net20
rlabel metal1 s 21418 4590 21418 4590 4 net21
rlabel metal1 s 18998 3026 18998 3026 4 net22
rlabel metal1 s 5520 2618 5520 2618 4 net23
rlabel metal1 s 14444 2550 14444 2550 4 net24
rlabel metal1 s 12708 5678 12708 5678 4 net25
rlabel metal1 s 4784 4182 4784 4182 4 net26
rlabel metal2 s 2639 7378 2639 7378 4 net27
rlabel metal2 s 2438 8738 2438 8738 4 net28
rlabel metal2 s 7406 11832 7406 11832 4 net29
rlabel metal1 s 2070 18394 2070 18394 4 net3
rlabel metal1 s 11638 2618 11638 2618 4 net30
rlabel metal2 s 10258 14280 10258 14280 4 net31
rlabel metal1 s 3749 12886 3749 12886 4 net32
rlabel metal2 s 4922 3910 4922 3910 4 net33
rlabel metal2 s 10350 7565 10350 7565 4 net34
rlabel metal2 s 2070 15912 2070 15912 4 net35
rlabel metal2 s 1903 18258 1903 18258 4 net36
rlabel metal1 s 4582 21522 4582 21522 4 net37
rlabel metal2 s 7774 22848 7774 22848 4 net38
rlabel metal1 s 10396 20570 10396 20570 4 net39
rlabel metal1 s 5336 21658 5336 21658 4 net4
rlabel metal1 s 10764 22950 10764 22950 4 net40
rlabel metal1 s 13276 16082 13276 16082 4 net41
rlabel metal1 s 13662 22984 13662 22984 4 net42
rlabel metal2 s 16496 22610 16496 22610 4 net43
rlabel metal1 s 19550 20910 19550 20910 4 net44
rlabel metal1 s 10028 2618 10028 2618 4 net45
rlabel metal2 s 21004 18258 21004 18258 4 net46
rlabel metal1 s 21068 15062 21068 15062 4 net47
rlabel metal1 s 21804 16422 21804 16422 4 net48
rlabel metal2 s 21850 13328 21850 13328 4 net49
rlabel metal2 s 8400 22610 8400 22610 4 net5
rlabel metal1 s 15134 11118 15134 11118 4 net50
rlabel metal2 s 19642 13022 19642 13022 4 net51
rlabel metal1 s 21188 10642 21188 10642 4 net52
rlabel metal1 s 21280 7378 21280 7378 4 net53
rlabel metal2 s 19440 3502 19440 3502 4 net54
rlabel metal1 s 17618 2618 17618 2618 4 net55
rlabel metal2 s 6946 2482 6946 2482 4 net56
rlabel metal2 s 14214 2924 14214 2924 4 net57
rlabel metal1 s 12880 2550 12880 2550 4 net58
rlabel metal1 s 4140 5542 4140 5542 4 net59
rlabel metal2 s 11086 21454 11086 21454 4 net6
rlabel metal2 s 1886 7480 1886 7480 4 net60
rlabel metal1 s 1748 10982 1748 10982 4 net61
rlabel metal1 s 7268 12818 7268 12818 4 net62
rlabel metal1 s 9246 2448 9246 2448 4 net63
rlabel metal1 s 10166 13226 10166 13226 4 net64
rlabel metal1 s 4048 12954 4048 12954 4 net65
rlabel metal2 s 4922 20978 4922 20978 4 net66
rlabel metal1 s 10350 2550 10350 2550 4 net67
rlabel metal2 s 5106 5746 5106 5746 4 net68
rlabel metal2 s 4922 19091 4922 19091 4 net69
rlabel metal1 s 11500 22950 11500 22950 4 net7
rlabel metal1 s 14122 2414 14122 2414 4 net70
rlabel metal1 s 16836 6154 16836 6154 4 net71
rlabel metal2 s 1702 8636 1702 8636 4 net72
rlabel metal1 s 5842 20978 5842 20978 4 net73
rlabel metal1 s 4922 18360 4922 18360 4 net74
rlabel metal1 s 6026 17238 6026 17238 4 net75
rlabel metal2 s 7222 19312 7222 19312 4 net76
rlabel metal1 s 7866 18394 7866 18394 4 net77
rlabel metal2 s 7038 18088 7038 18088 4 net78
rlabel metal2 s 17986 17867 17986 17867 4 net79
rlabel metal2 s 15364 17204 15364 17204 4 net8
rlabel metal1 s 13202 19482 13202 19482 4 net80
rlabel metal1 s 14214 23018 14214 23018 4 net81
rlabel metal2 s 16698 19363 16698 19363 4 net82
rlabel metal1 s 8556 2414 8556 2414 4 net83
rlabel metal1 s 16836 18122 16836 18122 4 net84
rlabel metal1 s 21252 18258 21252 18258 4 net85
rlabel metal2 s 21390 16830 21390 16830 4 net86
rlabel metal1 s 12190 15674 12190 15674 4 net87
rlabel metal1 s 15548 8330 15548 8330 4 net88
rlabel metal1 s 21298 6290 21298 6290 4 net89
rlabel metal1 s 13938 22032 13938 22032 4 net9
rlabel metal1 s 17894 9418 17894 9418 4 net90
rlabel metal1 s 21758 7922 21758 7922 4 net91
rlabel metal1 s 21390 8398 21390 8398 4 net92
rlabel metal1 s 15456 7174 15456 7174 4 net93
rlabel metal2 s 7866 4794 7866 4794 4 net94
rlabel metal1 s 16836 2414 16836 2414 4 net95
rlabel metal1 s 18952 8942 18952 8942 4 net96
rlabel metal2 s 3358 6154 3358 6154 4 net97
rlabel metal2 s 7452 4148 7452 4148 4 net98
rlabel metal1 s 1702 9996 1702 9996 4 net99
rlabel metal2 s 18722 1520 18722 1520 4 overflow
rlabel metal3 s 1096 8228 1096 8228 4 result[0]
rlabel metal3 s 1096 20468 1096 20468 4 result[10]
rlabel metal3 s 1096 17748 1096 17748 4 result[11]
rlabel metal3 s 0 17008 800 17128 4 result[12]
port 76 nsew
rlabel metal1 s 7268 23290 7268 23290 4 result[13]
rlabel metal2 s 8050 24123 8050 24123 4 result[14]
rlabel metal3 s 0 19728 800 19848 4 result[15]
port 79 nsew
rlabel metal2 s 18354 24123 18354 24123 4 result[16]
rlabel metal2 s 12282 24082 12282 24082 4 result[17]
rlabel metal1 s 14306 23290 14306 23290 4 result[18]
rlabel metal1 s 16560 23222 16560 23222 4 result[19]
rlabel metal2 s 8418 1520 8418 1520 4 result[1]
rlabel metal1 s 17112 23290 17112 23290 4 result[20]
rlabel metal2 s 21574 17901 21574 17901 4 result[21]
rlabel metal3 s 21574 17051 21574 17051 4 result[22]
rlabel metal2 s 11638 24116 11638 24116 4 result[23]
rlabel metal2 s 16146 1520 16146 1520 4 result[24]
rlabel metal3 s 21574 6171 21574 6171 4 result[25]
rlabel metal2 s 21942 9741 21942 9741 4 result[26]
rlabel metal2 s 21942 7633 21942 7633 4 result[27]
rlabel metal2 s 21574 8279 21574 8279 4 result[28]
rlabel metal2 s 15502 1520 15502 1520 4 result[29]
rlabel metal2 s 7774 1520 7774 1520 4 result[2]
rlabel metal2 s 16790 1520 16790 1520 4 result[30]
rlabel metal2 s 21942 8857 21942 8857 4 result[31]
rlabel metal3 s 1096 5508 1096 5508 4 result[3]
rlabel metal2 s 7130 1520 7130 1520 4 result[4]
rlabel metal3 s 1096 9588 1096 9588 4 result[5]
rlabel metal3 s 0 8848 800 8968 4 result[6]
port 101 nsew
rlabel metal2 s 5842 1520 5842 1520 4 result[7]
rlabel metal3 s 1096 19108 1096 19108 4 result[8]
rlabel metal3 s 0 15648 800 15768 4 result[9]
port 104 nsew
rlabel metal3 s 0 4088 800 4208 4 select[0]
port 105 nsew
rlabel metal3 s 0 21088 800 21208 4 select[1]
port 106 nsew
rlabel metal2 s 12926 1554 12926 1554 4 zero
flabel metal5 s 1056 21240 22404 21560 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 15936 22404 16256 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 10632 22404 10952 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 5328 22404 5648 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 20199 2128 20519 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 14886 2128 15206 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 9573 2128 9893 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4260 2128 4580 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 20580 22404 20900 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 15276 22404 15596 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 9972 22404 10292 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4668 22404 4988 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 19539 2128 19859 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 14226 2128 14546 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 8913 2128 9233 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3600 2128 3920 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 a[0]
port 3 nsew
flabel metal3 s 0 14968 800 15088 0 FreeSans 600 0 0 0 a[10]
port 4 nsew
flabel metal3 s 400 21828 400 21828 0 FreeSans 600 0 0 0 a[11]
flabel metal2 s 5170 24812 5226 25612 0 FreeSans 280 90 0 0 a[12]
port 6 nsew
flabel metal2 s 8390 24812 8446 25612 0 FreeSans 280 90 0 0 a[13]
port 7 nsew
flabel metal2 s 9034 24812 9090 25612 0 FreeSans 280 90 0 0 a[14]
port 8 nsew
flabel metal2 s 10966 24812 11022 25612 0 FreeSans 280 90 0 0 a[15]
port 9 nsew
flabel metal2 s 15474 24812 15530 25612 0 FreeSans 280 90 0 0 a[16]
port 10 nsew
flabel metal2 s 13542 24812 13598 25612 0 FreeSans 280 90 0 0 a[17]
port 11 nsew
flabel metal2 s 18694 24812 18750 25612 0 FreeSans 280 90 0 0 a[18]
port 12 nsew
flabel metal3 s 22668 20408 23468 20528 0 FreeSans 600 0 0 0 a[19]
port 13 nsew
flabel metal2 s 10966 0 11022 800 0 FreeSans 280 90 0 0 a[1]
port 14 nsew
flabel metal3 s 22668 19728 23468 19848 0 FreeSans 600 0 0 0 a[20]
port 15 nsew
flabel metal3 s 22668 15648 23468 15768 0 FreeSans 600 0 0 0 a[21]
port 16 nsew
flabel metal3 s 22668 19048 23468 19168 0 FreeSans 600 0 0 0 a[22]
port 17 nsew
flabel metal3 s 22668 12248 23468 12368 0 FreeSans 600 0 0 0 a[23]
port 18 nsew
flabel metal3 s 22668 11568 23468 11688 0 FreeSans 600 0 0 0 a[24]
port 19 nsew
flabel metal3 s 22668 14288 23468 14408 0 FreeSans 600 0 0 0 a[25]
port 20 nsew
flabel metal3 s 22668 4768 23468 4888 0 FreeSans 600 0 0 0 a[26]
port 21 nsew
flabel metal3 s 22668 5448 23468 5568 0 FreeSans 600 0 0 0 a[27]
port 22 nsew
flabel metal3 s 22668 4088 23468 4208 0 FreeSans 600 0 0 0 a[28]
port 23 nsew
flabel metal2 s 19982 0 20038 800 0 FreeSans 280 90 0 0 a[29]
port 24 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 a[2]
port 25 nsew
flabel metal2 s 17406 0 17462 800 0 FreeSans 280 90 0 0 a[30]
port 26 nsew
flabel metal2 s 12254 0 12310 800 0 FreeSans 280 90 0 0 a[31]
port 27 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 a[3]
port 28 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 a[4]
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 a[5]
flabel metal3 s 0 10888 800 11008 0 FreeSans 600 0 0 0 a[6]
port 31 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 a[7]
port 32 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 a[8]
port 33 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 a[9]
port 34 nsew
flabel metal3 s 400 3468 400 3468 0 FreeSans 600 0 0 0 ainv
flabel metal2 s 10322 0 10378 800 0 FreeSans 280 90 0 0 b[0]
port 36 nsew
flabel metal3 s 400 16388 400 16388 0 FreeSans 600 0 0 0 b[10]
flabel metal3 s 400 18428 400 18428 0 FreeSans 600 0 0 0 b[11]
flabel metal2 s 4526 24812 4582 25612 0 FreeSans 280 90 0 0 b[12]
port 39 nsew
flabel metal2 s 6458 24812 6514 25612 0 FreeSans 280 90 0 0 b[13]
port 40 nsew
flabel metal2 s 9678 24812 9734 25612 0 FreeSans 280 90 0 0 b[14]
port 41 nsew
flabel metal2 s 10322 24812 10378 25612 0 FreeSans 280 90 0 0 b[15]
port 42 nsew
flabel metal2 s 14830 24812 14886 25612 0 FreeSans 280 90 0 0 b[16]
port 43 nsew
flabel metal2 s 12898 24812 12954 25612 0 FreeSans 280 90 0 0 b[17]
port 44 nsew
flabel metal2 s 17406 24812 17462 25612 0 FreeSans 280 90 0 0 b[18]
port 45 nsew
flabel metal2 s 19338 24812 19394 25612 0 FreeSans 280 90 0 0 b[19]
port 46 nsew
flabel metal2 s 9678 0 9734 800 0 FreeSans 280 90 0 0 b[1]
port 47 nsew
flabel metal3 s 22668 18368 23468 18488 0 FreeSans 600 0 0 0 b[20]
port 48 nsew
flabel metal3 s 22668 14968 23468 15088 0 FreeSans 600 0 0 0 b[21]
port 49 nsew
flabel metal3 s 22668 16328 23468 16448 0 FreeSans 600 0 0 0 b[22]
port 50 nsew
flabel metal3 s 22668 13608 23468 13728 0 FreeSans 600 0 0 0 b[23]
port 51 nsew
flabel metal3 s 22668 10888 23468 11008 0 FreeSans 600 0 0 0 b[24]
port 52 nsew
flabel metal3 s 22668 12928 23468 13048 0 FreeSans 600 0 0 0 b[25]
port 53 nsew
flabel metal3 s 22668 10208 23468 10328 0 FreeSans 600 0 0 0 b[26]
port 54 nsew
flabel metal3 s 22668 6808 23468 6928 0 FreeSans 600 0 0 0 b[27]
port 55 nsew
flabel metal2 s 19338 0 19394 800 0 FreeSans 280 90 0 0 b[28]
port 56 nsew
flabel metal2 s 18050 0 18106 800 0 FreeSans 280 90 0 0 b[29]
port 57 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 b[2]
port 58 nsew
flabel metal2 s 14830 0 14886 800 0 FreeSans 280 90 0 0 b[30]
port 59 nsew
flabel metal2 s 13542 0 13598 800 0 FreeSans 280 90 0 0 b[31]
port 60 nsew
flabel metal3 s 400 4828 400 4828 0 FreeSans 600 0 0 0 b[3]
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 b[4]
port 62 nsew
flabel metal3 s 0 10208 800 10328 0 FreeSans 600 0 0 0 b[5]
port 63 nsew
flabel metal3 s 400 11628 400 11628 0 FreeSans 600 0 0 0 b[6]
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 b[7]
port 65 nsew
flabel metal3 s 400 14348 400 14348 0 FreeSans 600 0 0 0 b[8]
flabel metal3 s 400 12988 400 12988 0 FreeSans 600 0 0 0 b[9]
flabel metal3 s 400 22508 400 22508 0 FreeSans 600 0 0 0 binv
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 cin
port 69 nsew
flabel metal2 s 14186 0 14242 800 0 FreeSans 280 90 0 0 cout
port 70 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 fake_clk
port 71 nsew
flabel metal2 s 18694 0 18750 800 0 FreeSans 280 90 0 0 overflow
port 72 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 result[0]
port 73 nsew
flabel metal3 s 0 20408 800 20528 0 FreeSans 600 0 0 0 result[10]
port 74 nsew
flabel metal3 s 0 17688 800 17808 0 FreeSans 600 0 0 0 result[11]
port 75 nsew
flabel metal3 s 400 17068 400 17068 0 FreeSans 600 0 0 0 result[12]
flabel metal2 s 7102 24812 7158 25612 0 FreeSans 280 90 0 0 result[13]
port 77 nsew
flabel metal2 s 7746 24812 7802 25612 0 FreeSans 280 90 0 0 result[14]
port 78 nsew
flabel metal3 s 400 19788 400 19788 0 FreeSans 600 0 0 0 result[15]
flabel metal2 s 18050 24812 18106 25612 0 FreeSans 280 90 0 0 result[16]
port 80 nsew
flabel metal2 s 12254 24812 12310 25612 0 FreeSans 280 90 0 0 result[17]
port 81 nsew
flabel metal2 s 14186 24812 14242 25612 0 FreeSans 280 90 0 0 result[18]
port 82 nsew
flabel metal2 s 16118 24812 16174 25612 0 FreeSans 280 90 0 0 result[19]
port 83 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 result[1]
port 84 nsew
flabel metal2 s 16762 24812 16818 25612 0 FreeSans 280 90 0 0 result[20]
port 85 nsew
flabel metal3 s 22668 17688 23468 17808 0 FreeSans 600 0 0 0 result[21]
port 86 nsew
flabel metal3 s 22668 17008 23468 17128 0 FreeSans 600 0 0 0 result[22]
port 87 nsew
flabel metal2 s 11610 24812 11666 25612 0 FreeSans 280 90 0 0 result[23]
port 88 nsew
flabel metal2 s 16118 0 16174 800 0 FreeSans 280 90 0 0 result[24]
port 89 nsew
flabel metal3 s 22668 6128 23468 6248 0 FreeSans 600 0 0 0 result[25]
port 90 nsew
flabel metal3 s 22668 9528 23468 9648 0 FreeSans 600 0 0 0 result[26]
port 91 nsew
flabel metal3 s 22668 7488 23468 7608 0 FreeSans 600 0 0 0 result[27]
port 92 nsew
flabel metal3 s 22668 8168 23468 8288 0 FreeSans 600 0 0 0 result[28]
port 93 nsew
flabel metal2 s 15474 0 15530 800 0 FreeSans 280 90 0 0 result[29]
port 94 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 result[2]
port 95 nsew
flabel metal2 s 16762 0 16818 800 0 FreeSans 280 90 0 0 result[30]
port 96 nsew
flabel metal3 s 22668 8848 23468 8968 0 FreeSans 600 0 0 0 result[31]
port 97 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 result[3]
port 98 nsew
flabel metal2 s 7102 0 7158 800 0 FreeSans 280 90 0 0 result[4]
port 99 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 result[5]
port 100 nsew
flabel metal3 s 400 8908 400 8908 0 FreeSans 600 0 0 0 result[6]
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 result[7]
port 102 nsew
flabel metal3 s 0 19048 800 19168 0 FreeSans 600 0 0 0 result[8]
port 103 nsew
flabel metal3 s 400 15708 400 15708 0 FreeSans 600 0 0 0 result[9]
flabel metal3 s 400 4148 400 4148 0 FreeSans 600 0 0 0 select[0]
flabel metal3 s 400 21148 400 21148 0 FreeSans 600 0 0 0 select[1]
flabel metal2 s 12898 0 12954 800 0 FreeSans 280 90 0 0 zero
port 107 nsew
<< properties >>
string FIXED_BBOX 0 0 23468 25612
<< end >>
