magic
tech sky130A
magscale 1 2
timestamp 1743984720
<< checkpaint >>
rect -3932 -3932 29104 31248
<< viali >>
rect 5917 24769 5951 24803
rect 6561 24769 6595 24803
rect 7205 24769 7239 24803
rect 7849 24769 7883 24803
rect 8677 24769 8711 24803
rect 9321 24769 9355 24803
rect 9965 24769 9999 24803
rect 10609 24769 10643 24803
rect 11253 24769 11287 24803
rect 11713 24769 11747 24803
rect 12357 24769 12391 24803
rect 13001 24769 13035 24803
rect 13829 24769 13863 24803
rect 14473 24769 14507 24803
rect 15117 24769 15151 24803
rect 15761 24769 15795 24803
rect 16405 24769 16439 24803
rect 17049 24769 17083 24803
rect 17509 24769 17543 24803
rect 18153 24769 18187 24803
rect 20729 24769 20763 24803
rect 23673 24769 23707 24803
rect 22753 24701 22787 24735
rect 8493 24633 8527 24667
rect 9137 24633 9171 24667
rect 9781 24633 9815 24667
rect 10425 24633 10459 24667
rect 11069 24633 11103 24667
rect 14289 24633 14323 24667
rect 15577 24633 15611 24667
rect 16221 24633 16255 24667
rect 6101 24565 6135 24599
rect 6745 24565 6779 24599
rect 7389 24565 7423 24599
rect 8033 24565 8067 24599
rect 11897 24565 11931 24599
rect 12541 24565 12575 24599
rect 13185 24565 13219 24599
rect 13645 24565 13679 24599
rect 14933 24565 14967 24599
rect 16865 24565 16899 24599
rect 17693 24565 17727 24599
rect 18337 24565 18371 24599
rect 20913 24565 20947 24599
rect 23029 24225 23063 24259
rect 9070 24157 9104 24191
rect 14816 24157 14850 24191
rect 23673 24157 23707 24191
rect 8999 24021 9033 24055
rect 14887 24021 14921 24055
rect 8401 23817 8435 23851
rect 9321 23817 9355 23851
rect 14657 23817 14691 23851
rect 15577 23817 15611 23851
rect 17601 23817 17635 23851
rect 8493 23749 8527 23783
rect 15485 23749 15519 23783
rect 9413 23681 9447 23715
rect 9827 23681 9861 23715
rect 9930 23681 9964 23715
rect 17693 23681 17727 23715
rect 18107 23681 18141 23715
rect 18210 23681 18244 23715
rect 18454 23681 18488 23715
rect 23673 23681 23707 23715
rect 8309 23613 8343 23647
rect 9505 23613 9539 23647
rect 14749 23613 14783 23647
rect 14933 23613 14967 23647
rect 15669 23613 15703 23647
rect 17877 23613 17911 23647
rect 8861 23477 8895 23511
rect 8953 23477 8987 23511
rect 14289 23477 14323 23511
rect 15117 23477 15151 23511
rect 17233 23477 17267 23511
rect 18383 23477 18417 23511
rect 23489 23477 23523 23511
rect 14703 23273 14737 23307
rect 6929 23137 6963 23171
rect 17969 23137 18003 23171
rect 6745 23069 6779 23103
rect 7322 23069 7356 23103
rect 8953 23069 8987 23103
rect 9137 23069 9171 23103
rect 14806 23069 14840 23103
rect 17877 23069 17911 23103
rect 17785 23001 17819 23035
rect 6377 22933 6411 22967
rect 6837 22933 6871 22967
rect 7251 22933 7285 22967
rect 9321 22933 9355 22967
rect 17417 22933 17451 22967
rect 6929 22729 6963 22763
rect 7343 22729 7377 22763
rect 9505 22729 9539 22763
rect 12081 22729 12115 22763
rect 20453 22729 20487 22763
rect 14933 22661 14967 22695
rect 6837 22593 6871 22627
rect 7414 22593 7448 22627
rect 8585 22593 8619 22627
rect 9413 22593 9447 22627
rect 10057 22593 10091 22627
rect 12173 22593 12207 22627
rect 12587 22593 12621 22627
rect 12690 22593 12724 22627
rect 14473 22593 14507 22627
rect 15117 22593 15151 22627
rect 17233 22593 17267 22627
rect 20545 22593 20579 22627
rect 20959 22593 20993 22627
rect 21062 22593 21096 22627
rect 23673 22593 23707 22627
rect 7113 22525 7147 22559
rect 8677 22525 8711 22559
rect 9597 22525 9631 22559
rect 12357 22525 12391 22559
rect 14289 22525 14323 22559
rect 17049 22525 17083 22559
rect 20637 22525 20671 22559
rect 9873 22457 9907 22491
rect 6469 22389 6503 22423
rect 8953 22389 8987 22423
rect 9045 22389 9079 22423
rect 10241 22389 10275 22423
rect 11713 22389 11747 22423
rect 14657 22389 14691 22423
rect 14749 22389 14783 22423
rect 17417 22389 17451 22423
rect 20085 22389 20119 22423
rect 23489 22389 23523 22423
rect 9321 22185 9355 22219
rect 8953 22117 8987 22151
rect 9137 22049 9171 22083
rect 12633 22049 12667 22083
rect 14841 22049 14875 22083
rect 15025 22049 15059 22083
rect 15301 22049 15335 22083
rect 17509 22049 17543 22083
rect 17693 22049 17727 22083
rect 17969 22049 18003 22083
rect 12449 21981 12483 22015
rect 13026 21981 13060 22015
rect 14565 21981 14599 22015
rect 15393 21981 15427 22015
rect 16589 21981 16623 22015
rect 17233 21981 17267 22015
rect 18061 21981 18095 22015
rect 23673 21981 23707 22015
rect 6469 21913 6503 21947
rect 6653 21913 6687 21947
rect 16405 21913 16439 21947
rect 16773 21913 16807 21947
rect 17325 21913 17359 21947
rect 6837 21845 6871 21879
rect 12081 21845 12115 21879
rect 12541 21845 12575 21879
rect 12955 21845 12989 21879
rect 14197 21845 14231 21879
rect 14657 21845 14691 21879
rect 16865 21845 16899 21879
rect 23489 21845 23523 21879
rect 1593 21641 1627 21675
rect 3985 21573 4019 21607
rect 9873 21573 9907 21607
rect 1409 21505 1443 21539
rect 3376 21505 3410 21539
rect 3479 21505 3513 21539
rect 3893 21505 3927 21539
rect 4562 21505 4596 21539
rect 9137 21505 9171 21539
rect 9321 21505 9355 21539
rect 9689 21505 9723 21539
rect 12357 21505 12391 21539
rect 12541 21505 12575 21539
rect 14749 21505 14783 21539
rect 14933 21505 14967 21539
rect 15301 21505 15335 21539
rect 15485 21505 15519 21539
rect 17509 21505 17543 21539
rect 17693 21505 17727 21539
rect 17877 21505 17911 21539
rect 18061 21505 18095 21539
rect 18245 21505 18279 21539
rect 19625 21505 19659 21539
rect 23489 21505 23523 21539
rect 3801 21437 3835 21471
rect 6745 21437 6779 21471
rect 7205 21437 7239 21471
rect 11897 21437 11931 21471
rect 17325 21437 17359 21471
rect 19717 21437 19751 21471
rect 20085 21437 20119 21471
rect 20269 21437 20303 21471
rect 20729 21437 20763 21471
rect 20913 21437 20947 21471
rect 6561 21369 6595 21403
rect 7021 21369 7055 21403
rect 8953 21369 8987 21403
rect 12081 21369 12115 21403
rect 14565 21369 14599 21403
rect 20453 21369 20487 21403
rect 4353 21301 4387 21335
rect 4491 21301 4525 21335
rect 6929 21301 6963 21335
rect 7389 21301 7423 21335
rect 9505 21301 9539 21335
rect 11713 21301 11747 21335
rect 12173 21301 12207 21335
rect 15669 21301 15703 21335
rect 19993 21301 20027 21335
rect 20545 21301 20579 21335
rect 23673 21301 23707 21335
rect 15117 21097 15151 21131
rect 17785 21097 17819 21131
rect 10793 21029 10827 21063
rect 12725 21029 12759 21063
rect 21097 21029 21131 21063
rect 4445 20961 4479 20995
rect 4629 20961 4663 20995
rect 6101 20961 6135 20995
rect 6377 20961 6411 20995
rect 6929 20961 6963 20995
rect 7021 20961 7055 20995
rect 9229 20961 9263 20995
rect 9505 20961 9539 20995
rect 10425 20961 10459 20995
rect 10701 20961 10735 20995
rect 11253 20961 11287 20995
rect 11897 20961 11931 20995
rect 12081 20961 12115 20995
rect 12265 20961 12299 20995
rect 12909 20961 12943 20995
rect 14749 20961 14783 20995
rect 17049 20961 17083 20995
rect 17325 20961 17359 20995
rect 17417 20961 17451 20995
rect 17601 20961 17635 20995
rect 19073 20961 19107 20995
rect 19901 20961 19935 20995
rect 19993 20961 20027 20995
rect 20821 20961 20855 20995
rect 22753 20961 22787 20995
rect 1409 20893 1443 20927
rect 6009 20893 6043 20927
rect 7297 20893 7331 20927
rect 7665 20893 7699 20927
rect 9137 20893 9171 20927
rect 10333 20893 10367 20927
rect 11161 20893 11195 20927
rect 11805 20893 11839 20927
rect 12449 20893 12483 20927
rect 14933 20893 14967 20927
rect 16957 20893 16991 20927
rect 19809 20893 19843 20927
rect 21281 20893 21315 20927
rect 22477 20893 22511 20927
rect 23086 20893 23120 20927
rect 23673 20893 23707 20927
rect 4353 20825 4387 20859
rect 6837 20825 6871 20859
rect 7481 20825 7515 20859
rect 20637 20825 20671 20859
rect 21465 20825 21499 20859
rect 1593 20757 1627 20791
rect 3985 20757 4019 20791
rect 6469 20757 6503 20791
rect 11437 20757 11471 20791
rect 12633 20757 12667 20791
rect 13093 20757 13127 20791
rect 19441 20757 19475 20791
rect 20269 20757 20303 20791
rect 20729 20757 20763 20791
rect 22109 20757 22143 20791
rect 22569 20757 22603 20791
rect 22983 20757 23017 20791
rect 23489 20757 23523 20791
rect 6929 20553 6963 20587
rect 9137 20553 9171 20587
rect 14197 20553 14231 20587
rect 17233 20553 17267 20587
rect 19441 20553 19475 20587
rect 21005 20553 21039 20587
rect 12265 20485 12299 20519
rect 19349 20485 19383 20519
rect 20545 20485 20579 20519
rect 21373 20485 21407 20519
rect 3617 20417 3651 20451
rect 3801 20417 3835 20451
rect 4077 20417 4111 20451
rect 4537 20417 4571 20451
rect 6745 20417 6779 20451
rect 9229 20417 9263 20451
rect 9597 20417 9631 20451
rect 12081 20417 12115 20451
rect 15025 20417 15059 20451
rect 15117 20417 15151 20451
rect 15485 20417 15519 20451
rect 17325 20417 17359 20451
rect 17693 20417 17727 20451
rect 20269 20417 20303 20451
rect 20729 20417 20763 20451
rect 21189 20417 21223 20451
rect 4353 20349 4387 20383
rect 9413 20349 9447 20383
rect 14013 20349 14047 20383
rect 14105 20349 14139 20383
rect 15301 20349 15335 20383
rect 17509 20349 17543 20383
rect 19625 20349 19659 20383
rect 19901 20349 19935 20383
rect 20361 20349 20395 20383
rect 3893 20281 3927 20315
rect 6561 20281 6595 20315
rect 14657 20281 14691 20315
rect 3433 20213 3467 20247
rect 4261 20213 4295 20247
rect 4721 20213 4755 20247
rect 8769 20213 8803 20247
rect 10609 20213 10643 20247
rect 11897 20213 11931 20247
rect 14565 20213 14599 20247
rect 16865 20213 16899 20247
rect 18981 20213 19015 20247
rect 20913 20213 20947 20247
rect 14289 20009 14323 20043
rect 14933 20009 14967 20043
rect 16037 20009 16071 20043
rect 4169 19873 4203 19907
rect 6469 19873 6503 19907
rect 6929 19873 6963 19907
rect 9873 19873 9907 19907
rect 10609 19873 10643 19907
rect 10793 19873 10827 19907
rect 14657 19873 14691 19907
rect 16773 19873 16807 19907
rect 16957 19873 16991 19907
rect 1409 19805 1443 19839
rect 4353 19805 4387 19839
rect 4445 19805 4479 19839
rect 4905 19805 4939 19839
rect 5273 19805 5307 19839
rect 6561 19805 6595 19839
rect 7021 19805 7055 19839
rect 9689 19805 9723 19839
rect 14105 19805 14139 19839
rect 14565 19805 14599 19839
rect 15853 19805 15887 19839
rect 16681 19805 16715 19839
rect 23489 19805 23523 19839
rect 2605 19737 2639 19771
rect 5089 19737 5123 19771
rect 10517 19737 10551 19771
rect 4813 19669 4847 19703
rect 9321 19669 9355 19703
rect 9781 19669 9815 19703
rect 10149 19669 10183 19703
rect 16313 19669 16347 19703
rect 23673 19669 23707 19703
rect 7021 19465 7055 19499
rect 7113 19465 7147 19499
rect 8953 19465 8987 19499
rect 9045 19465 9079 19499
rect 18797 19465 18831 19499
rect 23397 19465 23431 19499
rect 23489 19465 23523 19499
rect 1593 19329 1627 19363
rect 3801 19329 3835 19363
rect 18613 19329 18647 19363
rect 23213 19329 23247 19363
rect 23673 19329 23707 19363
rect 3709 19261 3743 19295
rect 7297 19261 7331 19295
rect 8769 19261 8803 19295
rect 1409 19125 1443 19159
rect 4169 19125 4203 19159
rect 6653 19125 6687 19159
rect 9413 19125 9447 19159
rect 4169 18921 4203 18955
rect 7205 18921 7239 18955
rect 9137 18921 9171 18955
rect 9597 18921 9631 18955
rect 14381 18921 14415 18955
rect 18337 18921 18371 18955
rect 14657 18853 14691 18887
rect 3801 18785 3835 18819
rect 4445 18785 4479 18819
rect 6469 18785 6503 18819
rect 6653 18785 6687 18819
rect 12173 18785 12207 18819
rect 12357 18785 12391 18819
rect 12633 18785 12667 18819
rect 13001 18785 13035 18819
rect 13185 18785 13219 18819
rect 14289 18785 14323 18819
rect 14473 18785 14507 18819
rect 19809 18785 19843 18819
rect 21925 18785 21959 18819
rect 23213 18785 23247 18819
rect 1593 18717 1627 18751
rect 3985 18717 4019 18751
rect 4629 18717 4663 18751
rect 5089 18717 5123 18751
rect 6745 18717 6779 18751
rect 7389 18717 7423 18751
rect 8953 18717 8987 18751
rect 9413 18717 9447 18751
rect 11897 18717 11931 18751
rect 12725 18717 12759 18751
rect 17693 18717 17727 18751
rect 18153 18717 18187 18751
rect 20085 18717 20119 18751
rect 22937 18717 22971 18751
rect 23514 18717 23548 18751
rect 14105 18649 14139 18683
rect 14841 18649 14875 18683
rect 15025 18649 15059 18683
rect 19625 18649 19659 18683
rect 21741 18649 21775 18683
rect 1409 18581 1443 18615
rect 4537 18581 4571 18615
rect 4997 18581 5031 18615
rect 7113 18581 7147 18615
rect 11529 18581 11563 18615
rect 11989 18581 12023 18615
rect 13369 18581 13403 18615
rect 14197 18581 14231 18615
rect 19257 18581 19291 18615
rect 19717 18581 19751 18615
rect 21373 18581 21407 18615
rect 21833 18581 21867 18615
rect 22569 18581 22603 18615
rect 23029 18581 23063 18615
rect 23443 18581 23477 18615
rect 4261 18377 4295 18411
rect 4721 18377 4755 18411
rect 8861 18377 8895 18411
rect 14565 18377 14599 18411
rect 15301 18377 15335 18411
rect 17233 18377 17267 18411
rect 17785 18377 17819 18411
rect 18245 18377 18279 18411
rect 19533 18377 19567 18411
rect 19993 18377 20027 18411
rect 9505 18309 9539 18343
rect 13277 18309 13311 18343
rect 18153 18309 18187 18343
rect 22937 18309 22971 18343
rect 1593 18241 1627 18275
rect 3801 18241 3835 18275
rect 4629 18241 4663 18275
rect 9045 18241 9079 18275
rect 9229 18241 9263 18275
rect 11897 18241 11931 18275
rect 13093 18241 13127 18275
rect 14841 18241 14875 18275
rect 15761 18241 15795 18275
rect 15945 18241 15979 18275
rect 17325 18241 17359 18275
rect 19901 18241 19935 18275
rect 20729 18241 20763 18275
rect 22201 18241 22235 18275
rect 23029 18241 23063 18275
rect 23443 18241 23477 18275
rect 23546 18241 23580 18275
rect 3893 18173 3927 18207
rect 4169 18173 4203 18207
rect 4905 18173 4939 18207
rect 9137 18173 9171 18207
rect 14381 18173 14415 18207
rect 14749 18173 14783 18207
rect 15209 18173 15243 18207
rect 15485 18173 15519 18207
rect 17141 18173 17175 18207
rect 18337 18173 18371 18207
rect 20085 18173 20119 18207
rect 20361 18173 20395 18207
rect 20821 18173 20855 18207
rect 21005 18173 21039 18207
rect 21189 18173 21223 18207
rect 21833 18173 21867 18207
rect 22109 18173 22143 18207
rect 23121 18173 23155 18207
rect 9321 18105 9355 18139
rect 9505 18105 9539 18139
rect 13461 18105 13495 18139
rect 14197 18105 14231 18139
rect 15669 18105 15703 18139
rect 22569 18105 22603 18139
rect 1409 18037 1443 18071
rect 16129 18037 16163 18071
rect 17693 18037 17727 18071
rect 21373 18037 21407 18071
rect 6101 17833 6135 17867
rect 6561 17833 6595 17867
rect 9873 17833 9907 17867
rect 12633 17833 12667 17867
rect 13093 17833 13127 17867
rect 14749 17833 14783 17867
rect 16957 17833 16991 17867
rect 22109 17833 22143 17867
rect 22937 17833 22971 17867
rect 6837 17765 6871 17799
rect 9597 17765 9631 17799
rect 12725 17765 12759 17799
rect 21189 17765 21223 17799
rect 22477 17765 22511 17799
rect 23673 17765 23707 17799
rect 6377 17697 6411 17731
rect 7389 17697 7423 17731
rect 8217 17697 8251 17731
rect 10977 17697 11011 17731
rect 12357 17697 12391 17731
rect 15025 17697 15059 17731
rect 15669 17697 15703 17731
rect 16405 17697 16439 17731
rect 16497 17697 16531 17731
rect 22017 17697 22051 17731
rect 6285 17629 6319 17663
rect 6469 17629 6503 17663
rect 8125 17629 8159 17663
rect 8493 17629 8527 17663
rect 9413 17629 9447 17663
rect 9689 17629 9723 17663
rect 10885 17629 10919 17663
rect 12265 17629 12299 17663
rect 12909 17629 12943 17663
rect 15117 17629 15151 17663
rect 15853 17629 15887 17663
rect 17877 17629 17911 17663
rect 21373 17629 21407 17663
rect 21833 17629 21867 17663
rect 22293 17629 22327 17663
rect 22569 17629 22603 17663
rect 23489 17629 23523 17663
rect 6745 17561 6779 17595
rect 16037 17561 16071 17595
rect 16589 17561 16623 17595
rect 21557 17561 21591 17595
rect 21649 17561 21683 17595
rect 22753 17561 22787 17595
rect 6653 17493 6687 17527
rect 7205 17493 7239 17527
rect 7297 17493 7331 17527
rect 7665 17493 7699 17527
rect 8033 17493 8067 17527
rect 10425 17493 10459 17527
rect 10793 17493 10827 17527
rect 18061 17493 18095 17527
rect 5365 17289 5399 17323
rect 7021 17289 7055 17323
rect 11621 17289 11655 17323
rect 15117 17289 15151 17323
rect 15485 17221 15519 17255
rect 17969 17221 18003 17255
rect 1409 17153 1443 17187
rect 4997 17153 5031 17187
rect 7205 17153 7239 17187
rect 11989 17153 12023 17187
rect 12449 17153 12483 17187
rect 12633 17153 12667 17187
rect 13058 17153 13092 17187
rect 15577 17153 15611 17187
rect 15991 17153 16025 17187
rect 16094 17153 16128 17187
rect 16370 17145 16404 17179
rect 18061 17153 18095 17187
rect 18337 17153 18371 17187
rect 18889 17153 18923 17187
rect 23489 17153 23523 17187
rect 4813 17085 4847 17119
rect 4905 17085 4939 17119
rect 12081 17085 12115 17119
rect 12173 17085 12207 17119
rect 15761 17085 15795 17119
rect 18153 17085 18187 17119
rect 12817 17017 12851 17051
rect 19073 17017 19107 17051
rect 23673 17017 23707 17051
rect 1593 16949 1627 16983
rect 5457 16949 5491 16983
rect 12955 16949 12989 16983
rect 16267 16949 16301 16983
rect 18337 16949 18371 16983
rect 4813 16745 4847 16779
rect 7113 16745 7147 16779
rect 9413 16745 9447 16779
rect 11989 16745 12023 16779
rect 12449 16745 12483 16779
rect 15485 16745 15519 16779
rect 18429 16745 18463 16779
rect 19533 16745 19567 16779
rect 5273 16609 5307 16643
rect 5365 16609 5399 16643
rect 7757 16609 7791 16643
rect 9965 16609 9999 16643
rect 13093 16609 13127 16643
rect 15945 16609 15979 16643
rect 16037 16609 16071 16643
rect 17877 16609 17911 16643
rect 20085 16609 20119 16643
rect 1409 16541 1443 16575
rect 10241 16541 10275 16575
rect 12357 16541 12391 16575
rect 12817 16541 12851 16575
rect 13394 16541 13428 16575
rect 15853 16541 15887 16575
rect 18521 16541 18555 16575
rect 18797 16541 18831 16575
rect 20729 16541 20763 16575
rect 23673 16541 23707 16575
rect 9781 16473 9815 16507
rect 12173 16473 12207 16507
rect 1593 16405 1627 16439
rect 5181 16405 5215 16439
rect 7481 16405 7515 16439
rect 7573 16405 7607 16439
rect 9873 16405 9907 16439
rect 12909 16405 12943 16439
rect 13323 16405 13357 16439
rect 17969 16405 18003 16439
rect 18061 16405 18095 16439
rect 18705 16405 18739 16439
rect 19901 16405 19935 16439
rect 19993 16405 20027 16439
rect 23489 16405 23523 16439
rect 4353 16201 4387 16235
rect 7389 16201 7423 16235
rect 9689 16201 9723 16235
rect 10149 16201 10183 16235
rect 12357 16201 12391 16235
rect 12725 16201 12759 16235
rect 12817 16201 12851 16235
rect 14289 16201 14323 16235
rect 18153 16201 18187 16235
rect 18613 16201 18647 16235
rect 20361 16201 20395 16235
rect 20821 16201 20855 16235
rect 4169 16133 4203 16167
rect 1409 16065 1443 16099
rect 3985 16065 4019 16099
rect 4813 16065 4847 16099
rect 7021 16065 7055 16099
rect 7205 16065 7239 16099
rect 7665 16065 7699 16099
rect 10057 16065 10091 16099
rect 14105 16065 14139 16099
rect 18521 16065 18555 16099
rect 20729 16065 20763 16099
rect 22201 16065 22235 16099
rect 23673 16065 23707 16099
rect 4721 15997 4755 16031
rect 5181 15997 5215 16031
rect 7481 15997 7515 16031
rect 10333 15997 10367 16031
rect 13001 15997 13035 16031
rect 18705 15997 18739 16031
rect 20913 15997 20947 16031
rect 21833 15997 21867 16031
rect 22109 15997 22143 16031
rect 1593 15929 1627 15963
rect 7849 15861 7883 15895
rect 23489 15861 23523 15895
rect 3249 15657 3283 15691
rect 4997 15657 5031 15691
rect 5089 15657 5123 15691
rect 6929 15657 6963 15691
rect 7757 15657 7791 15691
rect 10057 15657 10091 15691
rect 14105 15657 14139 15691
rect 21005 15657 21039 15691
rect 1593 15589 1627 15623
rect 5457 15589 5491 15623
rect 6101 15589 6135 15623
rect 22201 15589 22235 15623
rect 3617 15521 3651 15555
rect 4445 15521 4479 15555
rect 6561 15521 6595 15555
rect 6745 15521 6779 15555
rect 7297 15521 7331 15555
rect 7573 15521 7607 15555
rect 8033 15521 8067 15555
rect 8585 15521 8619 15555
rect 8769 15521 8803 15555
rect 10701 15521 10735 15555
rect 14749 15521 14783 15555
rect 15577 15521 15611 15555
rect 18153 15521 18187 15555
rect 21557 15521 21591 15555
rect 1409 15453 1443 15487
rect 3433 15453 3467 15487
rect 5273 15453 5307 15487
rect 6285 15453 6319 15487
rect 7205 15453 7239 15487
rect 8125 15453 8159 15487
rect 15393 15453 15427 15487
rect 15761 15453 15795 15487
rect 17969 15453 18003 15487
rect 22017 15453 22051 15487
rect 23673 15453 23707 15487
rect 3801 15385 3835 15419
rect 3985 15385 4019 15419
rect 6469 15385 6503 15419
rect 8401 15385 8435 15419
rect 10425 15385 10459 15419
rect 4169 15317 4203 15351
rect 4537 15317 4571 15351
rect 4629 15317 4663 15351
rect 10517 15317 10551 15351
rect 14473 15317 14507 15351
rect 14565 15317 14599 15351
rect 14933 15317 14967 15351
rect 15301 15317 15335 15351
rect 17785 15317 17819 15351
rect 21373 15317 21407 15351
rect 21465 15317 21499 15351
rect 21833 15317 21867 15351
rect 23489 15317 23523 15351
rect 4721 15113 4755 15147
rect 7021 15113 7055 15147
rect 7389 15113 7423 15147
rect 9321 15113 9355 15147
rect 10609 15113 10643 15147
rect 10701 15113 10735 15147
rect 18429 15113 18463 15147
rect 20821 15113 20855 15147
rect 21465 15045 21499 15079
rect 22937 15045 22971 15079
rect 3893 14977 3927 15011
rect 9505 14977 9539 15011
rect 9689 14977 9723 15011
rect 9781 14977 9815 15011
rect 10241 14977 10275 15011
rect 10425 14977 10459 15011
rect 11932 14977 11966 15011
rect 18061 14977 18095 15011
rect 18889 14977 18923 15011
rect 21281 14977 21315 15011
rect 21649 14977 21683 15011
rect 22201 14977 22235 15011
rect 23029 14977 23063 15011
rect 23443 14977 23477 15011
rect 23546 14977 23580 15011
rect 3801 14909 3835 14943
rect 4261 14909 4295 14943
rect 4353 14909 4387 14943
rect 4537 14909 4571 14943
rect 7481 14909 7515 14943
rect 7665 14909 7699 14943
rect 9965 14909 9999 14943
rect 10885 14909 10919 14943
rect 17325 14909 17359 14943
rect 17785 14909 17819 14943
rect 17969 14909 18003 14943
rect 18521 14909 18555 14943
rect 18797 14909 18831 14943
rect 21005 14909 21039 14943
rect 21833 14909 21867 14943
rect 22109 14909 22143 14943
rect 23213 14909 23247 14943
rect 10149 14841 10183 14875
rect 11069 14841 11103 14875
rect 17509 14841 17543 14875
rect 21189 14841 21223 14875
rect 22569 14841 22603 14875
rect 12035 14773 12069 14807
rect 17141 14773 17175 14807
rect 3617 14569 3651 14603
rect 4261 14569 4295 14603
rect 6653 14569 6687 14603
rect 7527 14569 7561 14603
rect 9413 14569 9447 14603
rect 10517 14569 10551 14603
rect 11529 14569 11563 14603
rect 12357 14569 12391 14603
rect 14841 14569 14875 14603
rect 15117 14569 15151 14603
rect 17969 14569 18003 14603
rect 18429 14569 18463 14603
rect 21465 14569 21499 14603
rect 21925 14569 21959 14603
rect 9873 14501 9907 14535
rect 22293 14501 22327 14535
rect 3065 14433 3099 14467
rect 4905 14433 4939 14467
rect 7205 14433 7239 14467
rect 9597 14433 9631 14467
rect 9781 14433 9815 14467
rect 10333 14433 10367 14467
rect 10793 14433 10827 14467
rect 12173 14433 12207 14467
rect 12817 14433 12851 14467
rect 13001 14433 13035 14467
rect 14197 14433 14231 14467
rect 15577 14433 15611 14467
rect 17693 14433 17727 14467
rect 19901 14433 19935 14467
rect 23121 14433 23155 14467
rect 1409 14365 1443 14399
rect 3249 14365 3283 14399
rect 3934 14365 3968 14399
rect 5206 14365 5240 14399
rect 7021 14365 7055 14399
rect 7598 14365 7632 14399
rect 7874 14365 7908 14399
rect 10241 14365 10275 14399
rect 10885 14365 10919 14399
rect 13553 14365 13587 14399
rect 15485 14365 15519 14399
rect 16957 14365 16991 14399
rect 17141 14365 17175 14399
rect 17325 14365 17359 14399
rect 17601 14365 17635 14399
rect 18061 14365 18095 14399
rect 18940 14365 18974 14399
rect 19625 14365 19659 14399
rect 21649 14365 21683 14399
rect 22109 14365 22143 14399
rect 22937 14365 22971 14399
rect 23514 14365 23548 14399
rect 3157 14297 3191 14331
rect 3847 14297 3881 14331
rect 12725 14297 12759 14331
rect 13737 14297 13771 14331
rect 18245 14297 18279 14331
rect 19027 14297 19061 14331
rect 19717 14297 19751 14331
rect 21833 14297 21867 14331
rect 1593 14229 1627 14263
rect 4629 14229 4663 14263
rect 4721 14229 4755 14263
rect 5135 14229 5169 14263
rect 7113 14229 7147 14263
rect 7803 14229 7837 14263
rect 11897 14229 11931 14263
rect 11989 14229 12023 14263
rect 13921 14229 13955 14263
rect 14381 14229 14415 14263
rect 14473 14229 14507 14263
rect 19257 14229 19291 14263
rect 22569 14229 22603 14263
rect 23029 14229 23063 14263
rect 23443 14229 23477 14263
rect 1593 14025 1627 14059
rect 11943 14025 11977 14059
rect 14197 14025 14231 14059
rect 17601 14025 17635 14059
rect 18061 14025 18095 14059
rect 1409 13889 1443 13923
rect 12014 13889 12048 13923
rect 14473 13889 14507 13923
rect 15485 13889 15519 13923
rect 17233 13889 17267 13923
rect 17877 13889 17911 13923
rect 23397 13889 23431 13923
rect 23673 13889 23707 13923
rect 13829 13821 13863 13855
rect 14013 13821 14047 13855
rect 14381 13821 14415 13855
rect 14841 13821 14875 13855
rect 15669 13821 15703 13855
rect 17049 13821 17083 13855
rect 17141 13821 17175 13855
rect 17693 13821 17727 13855
rect 23489 13753 23523 13787
rect 15301 13685 15335 13719
rect 23213 13685 23247 13719
rect 13829 13481 13863 13515
rect 17187 13481 17221 13515
rect 14381 13413 14415 13447
rect 23489 13413 23523 13447
rect 13185 13345 13219 13379
rect 14565 13345 14599 13379
rect 19625 13345 19659 13379
rect 1409 13277 1443 13311
rect 6996 13277 7030 13311
rect 13461 13277 13495 13311
rect 14254 13277 14288 13311
rect 15485 13277 15519 13311
rect 17258 13277 17292 13311
rect 19441 13277 19475 13311
rect 20970 13277 21004 13311
rect 23673 13277 23707 13311
rect 13369 13209 13403 13243
rect 14151 13209 14185 13243
rect 14749 13209 14783 13243
rect 15301 13209 15335 13243
rect 1593 13141 1627 13175
rect 7067 13141 7101 13175
rect 15669 13141 15703 13175
rect 19257 13141 19291 13175
rect 20867 13141 20901 13175
rect 6929 12937 6963 12971
rect 10241 12937 10275 12971
rect 14381 12937 14415 12971
rect 19165 12937 19199 12971
rect 20269 12937 20303 12971
rect 20637 12937 20671 12971
rect 20729 12937 20763 12971
rect 8493 12869 8527 12903
rect 19809 12869 19843 12903
rect 19993 12869 20027 12903
rect 1409 12801 1443 12835
rect 4420 12801 4454 12835
rect 4997 12801 5031 12835
rect 5089 12801 5123 12835
rect 5503 12801 5537 12835
rect 5606 12801 5640 12835
rect 7021 12801 7055 12835
rect 8585 12801 8619 12835
rect 8999 12801 9033 12835
rect 9102 12801 9136 12835
rect 10425 12801 10459 12835
rect 10609 12801 10643 12835
rect 14013 12801 14047 12835
rect 14622 12801 14656 12835
rect 19257 12801 19291 12835
rect 19625 12801 19659 12835
rect 21246 12801 21280 12835
rect 23673 12801 23707 12835
rect 5273 12733 5307 12767
rect 6837 12733 6871 12767
rect 7849 12733 7883 12767
rect 8677 12733 8711 12767
rect 13829 12733 13863 12767
rect 13921 12733 13955 12767
rect 14519 12733 14553 12767
rect 19349 12733 19383 12767
rect 20821 12733 20855 12767
rect 1593 12665 1627 12699
rect 4491 12665 4525 12699
rect 7389 12665 7423 12699
rect 7665 12665 7699 12699
rect 8033 12665 8067 12699
rect 23489 12665 23523 12699
rect 4629 12597 4663 12631
rect 8125 12597 8159 12631
rect 18797 12597 18831 12631
rect 21143 12597 21177 12631
rect 9689 12393 9723 12427
rect 6837 12325 6871 12359
rect 10793 12325 10827 12359
rect 19901 12325 19935 12359
rect 4629 12257 4663 12291
rect 4721 12257 4755 12291
rect 8033 12257 8067 12291
rect 8677 12257 8711 12291
rect 9321 12257 9355 12291
rect 10057 12257 10091 12291
rect 10333 12257 10367 12291
rect 11253 12257 11287 12291
rect 15669 12257 15703 12291
rect 16037 12257 16071 12291
rect 19257 12257 19291 12291
rect 19533 12257 19567 12291
rect 20913 12257 20947 12291
rect 21097 12257 21131 12291
rect 6653 12189 6687 12223
rect 6929 12189 6963 12223
rect 7113 12189 7147 12223
rect 7297 12189 7331 12223
rect 7849 12189 7883 12223
rect 8309 12189 8343 12223
rect 9505 12189 9539 12223
rect 9965 12189 9999 12223
rect 10425 12189 10459 12223
rect 11161 12189 11195 12223
rect 12506 12189 12540 12223
rect 15853 12189 15887 12223
rect 16380 12189 16414 12223
rect 19625 12189 19659 12223
rect 20085 12189 20119 12223
rect 20821 12189 20855 12223
rect 7757 12121 7791 12155
rect 8493 12121 8527 12155
rect 11621 12121 11655 12155
rect 11805 12121 11839 12155
rect 4813 12053 4847 12087
rect 5181 12053 5215 12087
rect 6469 12053 6503 12087
rect 7389 12053 7423 12087
rect 11437 12053 11471 12087
rect 12403 12053 12437 12087
rect 16451 12053 16485 12087
rect 20269 12053 20303 12087
rect 20453 12053 20487 12087
rect 1593 11849 1627 11883
rect 8309 11849 8343 11883
rect 10241 11849 10275 11883
rect 10333 11849 10367 11883
rect 10885 11849 10919 11883
rect 17141 11849 17175 11883
rect 23489 11849 23523 11883
rect 3801 11781 3835 11815
rect 5089 11781 5123 11815
rect 12541 11781 12575 11815
rect 17049 11781 17083 11815
rect 20177 11781 20211 11815
rect 1409 11713 1443 11747
rect 3985 11713 4019 11747
rect 4261 11713 4295 11747
rect 4445 11713 4479 11747
rect 5733 11713 5767 11747
rect 7481 11713 7515 11747
rect 12633 11713 12667 11747
rect 13047 11713 13081 11747
rect 13150 11713 13184 11747
rect 15577 11713 15611 11747
rect 18521 11713 18555 11747
rect 18981 11713 19015 11747
rect 19165 11713 19199 11747
rect 19993 11713 20027 11747
rect 23673 11713 23707 11747
rect 4629 11645 4663 11679
rect 5181 11645 5215 11679
rect 5365 11645 5399 11679
rect 5549 11645 5583 11679
rect 7389 11645 7423 11679
rect 8125 11645 8159 11679
rect 10517 11645 10551 11679
rect 11069 11645 11103 11679
rect 11713 11645 11747 11679
rect 12817 11645 12851 11679
rect 15669 11645 15703 11679
rect 16221 11645 16255 11679
rect 17233 11645 17267 11679
rect 18613 11645 18647 11679
rect 4169 11577 4203 11611
rect 7941 11577 7975 11611
rect 11253 11577 11287 11611
rect 11897 11577 11931 11611
rect 12173 11577 12207 11611
rect 16037 11577 16071 11611
rect 16681 11577 16715 11611
rect 18797 11577 18831 11611
rect 4721 11509 4755 11543
rect 5917 11509 5951 11543
rect 7849 11509 7883 11543
rect 9873 11509 9907 11543
rect 11529 11509 11563 11543
rect 15945 11509 15979 11543
rect 16405 11509 16439 11543
rect 18153 11509 18187 11543
rect 19809 11509 19843 11543
rect 1593 11305 1627 11339
rect 11989 11305 12023 11339
rect 14933 11305 14967 11339
rect 16865 11305 16899 11339
rect 9597 11237 9631 11271
rect 11161 11237 11195 11271
rect 23489 11237 23523 11271
rect 4813 11169 4847 11203
rect 5089 11169 5123 11203
rect 5457 11169 5491 11203
rect 7665 11169 7699 11203
rect 7941 11169 7975 11203
rect 10057 11169 10091 11203
rect 10149 11169 10183 11203
rect 11621 11169 11655 11203
rect 11713 11169 11747 11203
rect 12449 11169 12483 11203
rect 12633 11169 12667 11203
rect 14289 11169 14323 11203
rect 15945 11169 15979 11203
rect 16221 11169 16255 11203
rect 18429 11169 18463 11203
rect 22109 11169 22143 11203
rect 1409 11101 1443 11135
rect 4721 11101 4755 11135
rect 5825 11101 5859 11135
rect 7573 11101 7607 11135
rect 9965 11101 9999 11135
rect 11529 11101 11563 11135
rect 14565 11101 14599 11135
rect 15163 11101 15197 11135
rect 15853 11101 15887 11135
rect 16681 11101 16715 11135
rect 18245 11101 18279 11135
rect 18705 11101 18739 11135
rect 21925 11101 21959 11135
rect 22994 11101 23028 11135
rect 23673 11101 23707 11135
rect 5641 11033 5675 11067
rect 12357 11033 12391 11067
rect 14473 11033 14507 11067
rect 15071 11033 15105 11067
rect 16497 11033 16531 11067
rect 21281 11033 21315 11067
rect 21465 11033 21499 11067
rect 21649 11033 21683 11067
rect 21741 11033 21775 11067
rect 17877 10965 17911 10999
rect 18337 10965 18371 10999
rect 22891 10965 22925 10999
rect 5825 10761 5859 10795
rect 13369 10761 13403 10795
rect 13829 10761 13863 10795
rect 14013 10761 14047 10795
rect 18061 10761 18095 10795
rect 18429 10761 18463 10795
rect 18521 10761 18555 10795
rect 15301 10693 15335 10727
rect 15485 10693 15519 10727
rect 23029 10693 23063 10727
rect 1593 10625 1627 10659
rect 4997 10625 5031 10659
rect 13185 10625 13219 10659
rect 13277 10625 13311 10659
rect 13645 10625 13679 10659
rect 13737 10625 13771 10659
rect 14013 10625 14047 10659
rect 14105 10625 14139 10659
rect 14289 10625 14323 10659
rect 15945 10625 15979 10659
rect 20729 10625 20763 10659
rect 21465 10625 21499 10659
rect 22201 10625 22235 10659
rect 23121 10625 23155 10659
rect 23535 10625 23569 10659
rect 23638 10625 23672 10659
rect 5089 10557 5123 10591
rect 5641 10557 5675 10591
rect 13553 10557 13587 10591
rect 15761 10557 15795 10591
rect 18705 10557 18739 10591
rect 20821 10557 20855 10591
rect 21097 10557 21131 10591
rect 21557 10557 21591 10591
rect 22293 10557 22327 10591
rect 22385 10557 22419 10591
rect 23213 10557 23247 10591
rect 5457 10489 5491 10523
rect 13461 10489 13495 10523
rect 21833 10489 21867 10523
rect 1409 10421 1443 10455
rect 5365 10421 5399 10455
rect 14289 10421 14323 10455
rect 15669 10421 15703 10455
rect 16129 10421 16163 10455
rect 19993 10421 20027 10455
rect 20361 10421 20395 10455
rect 22661 10421 22695 10455
rect 21281 10217 21315 10251
rect 22017 10217 22051 10251
rect 22109 10217 22143 10251
rect 23489 10217 23523 10251
rect 5457 10081 5491 10115
rect 6837 10081 6871 10115
rect 8125 10081 8159 10115
rect 15853 10081 15887 10115
rect 16037 10081 16071 10115
rect 19809 10081 19843 10115
rect 20545 10081 20579 10115
rect 20637 10081 20671 10115
rect 20913 10081 20947 10115
rect 21097 10081 21131 10115
rect 22477 10081 22511 10115
rect 23029 10081 23063 10115
rect 23121 10081 23155 10115
rect 1593 10013 1627 10047
rect 5273 10013 5307 10047
rect 5365 10013 5399 10047
rect 5733 10013 5767 10047
rect 7021 10013 7055 10047
rect 7849 10013 7883 10047
rect 7941 10013 7975 10047
rect 8309 10013 8343 10047
rect 15761 10013 15795 10047
rect 17693 10013 17727 10047
rect 19625 10013 19659 10047
rect 20453 10013 20487 10047
rect 21649 10013 21683 10047
rect 22293 10013 22327 10047
rect 23673 10013 23707 10047
rect 6929 9945 6963 9979
rect 21833 9945 21867 9979
rect 1409 9877 1443 9911
rect 4905 9877 4939 9911
rect 7389 9877 7423 9911
rect 7481 9877 7515 9911
rect 15393 9877 15427 9911
rect 17877 9877 17911 9911
rect 19257 9877 19291 9911
rect 19717 9877 19751 9911
rect 20085 9877 20119 9911
rect 22569 9877 22603 9911
rect 22937 9877 22971 9911
rect 4905 9673 4939 9707
rect 7481 9673 7515 9707
rect 15669 9673 15703 9707
rect 17325 9673 17359 9707
rect 4997 9605 5031 9639
rect 7021 9605 7055 9639
rect 17601 9605 17635 9639
rect 5641 9537 5675 9571
rect 7665 9537 7699 9571
rect 10425 9537 10459 9571
rect 11002 9537 11036 9571
rect 13461 9537 13495 9571
rect 16681 9537 16715 9571
rect 17233 9537 17267 9571
rect 17509 9537 17543 9571
rect 17969 9537 18003 9571
rect 23489 9537 23523 9571
rect 4813 9469 4847 9503
rect 7205 9469 7239 9503
rect 7389 9469 7423 9503
rect 9781 9469 9815 9503
rect 9965 9469 9999 9503
rect 10517 9469 10551 9503
rect 13277 9469 13311 9503
rect 13369 9469 13403 9503
rect 15485 9469 15519 9503
rect 15577 9469 15611 9503
rect 5365 9401 5399 9435
rect 7021 9401 7055 9435
rect 10793 9401 10827 9435
rect 13829 9401 13863 9435
rect 18153 9401 18187 9435
rect 23673 9401 23707 9435
rect 5457 9333 5491 9367
rect 7297 9333 7331 9367
rect 9597 9333 9631 9367
rect 10931 9333 10965 9367
rect 13921 9333 13955 9367
rect 16037 9333 16071 9367
rect 16221 9333 16255 9367
rect 16865 9333 16899 9367
rect 17417 9333 17451 9367
rect 8033 9129 8067 9163
rect 13737 9129 13771 9163
rect 15761 9129 15795 9163
rect 1409 9061 1443 9095
rect 7757 9061 7791 9095
rect 11621 9061 11655 9095
rect 17785 9061 17819 9095
rect 8493 8993 8527 9027
rect 8585 8993 8619 9027
rect 9781 8993 9815 9027
rect 11069 8993 11103 9027
rect 12173 8993 12207 9027
rect 13185 8993 13219 9027
rect 13277 8993 13311 9027
rect 16221 8993 16255 9027
rect 16405 8993 16439 9027
rect 1593 8925 1627 8959
rect 7941 8925 7975 8959
rect 9505 8925 9539 8959
rect 11370 8925 11404 8959
rect 17601 8925 17635 8959
rect 23489 8925 23523 8959
rect 8401 8857 8435 8891
rect 10149 8857 10183 8891
rect 10333 8857 10367 8891
rect 10793 8857 10827 8891
rect 16129 8857 16163 8891
rect 9137 8789 9171 8823
rect 9597 8789 9631 8823
rect 9965 8789 9999 8823
rect 10425 8789 10459 8823
rect 10885 8789 10919 8823
rect 11299 8789 11333 8823
rect 11989 8789 12023 8823
rect 12081 8789 12115 8823
rect 13369 8789 13403 8823
rect 23673 8789 23707 8823
rect 5273 8585 5307 8619
rect 10793 8585 10827 8619
rect 13185 8585 13219 8619
rect 17877 8585 17911 8619
rect 18337 8585 18371 8619
rect 18705 8585 18739 8619
rect 4721 8449 4755 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 10057 8449 10091 8483
rect 10241 8449 10275 8483
rect 10701 8449 10735 8483
rect 11713 8449 11747 8483
rect 13553 8449 13587 8483
rect 15577 8449 15611 8483
rect 16681 8449 16715 8483
rect 18245 8449 18279 8483
rect 19073 8449 19107 8483
rect 19165 8449 19199 8483
rect 19533 8449 19567 8483
rect 22017 8449 22051 8483
rect 22201 8449 22235 8483
rect 22962 8449 22996 8483
rect 23489 8449 23523 8483
rect 4537 8381 4571 8415
rect 10977 8381 11011 8415
rect 11621 8381 11655 8415
rect 12081 8381 12115 8415
rect 13645 8381 13679 8415
rect 13737 8381 13771 8415
rect 18521 8381 18555 8415
rect 19257 8381 19291 8415
rect 22477 8381 22511 8415
rect 22661 8381 22695 8415
rect 4353 8313 4387 8347
rect 9873 8313 9907 8347
rect 15761 8313 15795 8347
rect 23673 8313 23707 8347
rect 10333 8245 10367 8279
rect 16865 8245 16899 8279
rect 20913 8245 20947 8279
rect 21833 8245 21867 8279
rect 22293 8245 22327 8279
rect 22891 8245 22925 8279
rect 5641 8041 5675 8075
rect 10149 8041 10183 8075
rect 13461 8041 13495 8075
rect 13921 8041 13955 8075
rect 15393 8041 15427 8075
rect 19533 8041 19567 8075
rect 22569 8041 22603 8075
rect 10885 7973 10919 8007
rect 4445 7905 4479 7939
rect 4721 7905 4755 7939
rect 4997 7905 5031 7939
rect 6009 7905 6043 7939
rect 10517 7905 10551 7939
rect 11069 7905 11103 7939
rect 11253 7905 11287 7939
rect 13553 7905 13587 7939
rect 14657 7905 14691 7939
rect 15577 7905 15611 7939
rect 15761 7905 15795 7939
rect 20085 7905 20119 7939
rect 20913 7905 20947 7939
rect 21097 7905 21131 7939
rect 21741 7905 21775 7939
rect 21833 7905 21867 7939
rect 22109 7905 22143 7939
rect 23121 7905 23155 7939
rect 1409 7837 1443 7871
rect 4353 7837 4387 7871
rect 5825 7837 5859 7871
rect 7205 7837 7239 7871
rect 10333 7837 10367 7871
rect 13093 7837 13127 7871
rect 13737 7837 13771 7871
rect 15669 7837 15703 7871
rect 22293 7837 22327 7871
rect 22937 7837 22971 7871
rect 23514 7837 23548 7871
rect 13277 7769 13311 7803
rect 14473 7769 14507 7803
rect 15393 7769 15427 7803
rect 19901 7769 19935 7803
rect 1593 7701 1627 7735
rect 5089 7701 5123 7735
rect 5181 7701 5215 7735
rect 5549 7701 5583 7735
rect 14105 7701 14139 7735
rect 14565 7701 14599 7735
rect 19993 7701 20027 7735
rect 20453 7701 20487 7735
rect 20821 7701 20855 7735
rect 21281 7701 21315 7735
rect 21649 7701 21683 7735
rect 22477 7701 22511 7735
rect 23029 7701 23063 7735
rect 23443 7701 23477 7735
rect 1593 7497 1627 7531
rect 3709 7497 3743 7531
rect 5365 7497 5399 7531
rect 7297 7497 7331 7531
rect 9045 7497 9079 7531
rect 14059 7497 14093 7531
rect 22569 7497 22603 7531
rect 22937 7497 22971 7531
rect 23029 7497 23063 7531
rect 23489 7497 23523 7531
rect 3341 7429 3375 7463
rect 4537 7429 4571 7463
rect 4997 7429 5031 7463
rect 1409 7361 1443 7395
rect 2732 7361 2766 7395
rect 2835 7361 2869 7395
rect 3249 7361 3283 7395
rect 3928 7361 3962 7395
rect 4031 7361 4065 7395
rect 4445 7361 4479 7395
rect 5181 7361 5215 7395
rect 5825 7361 5859 7395
rect 7205 7361 7239 7395
rect 7849 7361 7883 7395
rect 9137 7361 9171 7395
rect 9413 7361 9447 7395
rect 13988 7361 14022 7395
rect 15301 7361 15335 7395
rect 15945 7361 15979 7395
rect 18705 7361 18739 7395
rect 21465 7361 21499 7395
rect 22201 7361 22235 7395
rect 23673 7361 23707 7395
rect 3157 7293 3191 7327
rect 4261 7293 4295 7327
rect 5733 7293 5767 7327
rect 6193 7293 6227 7327
rect 7389 7293 7423 7327
rect 8769 7293 8803 7327
rect 8953 7293 8987 7327
rect 18797 7293 18831 7327
rect 19073 7293 19107 7327
rect 21097 7293 21131 7327
rect 21557 7293 21591 7327
rect 21833 7293 21867 7327
rect 22109 7293 22143 7327
rect 23213 7293 23247 7327
rect 4905 7225 4939 7259
rect 15485 7225 15519 7259
rect 6837 7157 6871 7191
rect 8033 7157 8067 7191
rect 8861 7157 8895 7191
rect 9229 7157 9263 7191
rect 16129 7157 16163 7191
rect 4813 6953 4847 6987
rect 7481 6953 7515 6987
rect 16313 6953 16347 6987
rect 4445 6885 4479 6919
rect 13737 6885 13771 6919
rect 22201 6885 22235 6919
rect 4629 6817 4663 6851
rect 6929 6817 6963 6851
rect 13001 6817 13035 6851
rect 13277 6817 13311 6851
rect 15669 6817 15703 6851
rect 16957 6817 16991 6851
rect 17785 6817 17819 6851
rect 19073 6817 19107 6851
rect 21373 6817 21407 6851
rect 22017 6817 22051 6851
rect 7021 6749 7055 6783
rect 7113 6749 7147 6783
rect 7757 6749 7791 6783
rect 8401 6749 8435 6783
rect 9597 6749 9631 6783
rect 10885 6749 10919 6783
rect 12909 6749 12943 6783
rect 13553 6749 13587 6783
rect 17601 6749 17635 6783
rect 17969 6749 18003 6783
rect 18889 6749 18923 6783
rect 21557 6749 21591 6783
rect 23489 6749 23523 6783
rect 15393 6681 15427 6715
rect 21741 6681 21775 6715
rect 21833 6681 21867 6715
rect 7573 6613 7607 6647
rect 8585 6613 8619 6647
rect 9781 6613 9815 6647
rect 13369 6613 13403 6647
rect 15025 6613 15059 6647
rect 15485 6613 15519 6647
rect 16681 6613 16715 6647
rect 16773 6613 16807 6647
rect 17141 6613 17175 6647
rect 17509 6613 17543 6647
rect 18705 6613 18739 6647
rect 23673 6613 23707 6647
rect 8125 6409 8159 6443
rect 8677 6409 8711 6443
rect 9689 6409 9723 6443
rect 10149 6409 10183 6443
rect 10517 6409 10551 6443
rect 10977 6409 11011 6443
rect 13185 6409 13219 6443
rect 15393 6409 15427 6443
rect 18797 6409 18831 6443
rect 23489 6409 23523 6443
rect 12817 6341 12851 6375
rect 18521 6341 18555 6375
rect 8217 6273 8251 6307
rect 9045 6273 9079 6307
rect 10057 6273 10091 6307
rect 10885 6273 10919 6307
rect 13645 6273 13679 6307
rect 14105 6273 14139 6307
rect 15761 6273 15795 6307
rect 15853 6273 15887 6307
rect 16221 6273 16255 6307
rect 18705 6273 18739 6307
rect 19165 6273 19199 6307
rect 19993 6273 20027 6307
rect 23673 6273 23707 6307
rect 7941 6205 7975 6239
rect 9137 6205 9171 6239
rect 9229 6205 9263 6239
rect 10241 6205 10275 6239
rect 11069 6205 11103 6239
rect 12541 6205 12575 6239
rect 12725 6205 12759 6239
rect 13553 6205 13587 6239
rect 14197 6205 14231 6239
rect 16037 6205 16071 6239
rect 19257 6205 19291 6239
rect 19349 6205 19383 6239
rect 20085 6205 20119 6239
rect 8585 6137 8619 6171
rect 19625 6137 19659 6171
rect 13277 6069 13311 6103
rect 14473 6069 14507 6103
rect 18337 6069 18371 6103
rect 5549 5865 5583 5899
rect 8677 5865 8711 5899
rect 11069 5865 11103 5899
rect 12771 5865 12805 5899
rect 17233 5865 17267 5899
rect 18705 5865 18739 5899
rect 19717 5865 19751 5899
rect 23489 5865 23523 5899
rect 11161 5797 11195 5831
rect 4997 5729 5031 5763
rect 10793 5729 10827 5763
rect 13737 5729 13771 5763
rect 13921 5729 13955 5763
rect 17693 5729 17727 5763
rect 19073 5729 19107 5763
rect 19257 5729 19291 5763
rect 19625 5729 19659 5763
rect 5641 5661 5675 5695
rect 10701 5661 10735 5695
rect 11345 5661 11379 5695
rect 12874 5661 12908 5695
rect 13461 5661 13495 5695
rect 17601 5661 17635 5695
rect 18889 5661 18923 5695
rect 19441 5661 19475 5695
rect 20085 5661 20119 5695
rect 23673 5661 23707 5695
rect 13277 5593 13311 5627
rect 13553 5593 13587 5627
rect 19901 5593 19935 5627
rect 5089 5525 5123 5559
rect 5181 5525 5215 5559
rect 11529 5525 11563 5559
rect 13093 5525 13127 5559
rect 5089 5321 5123 5355
rect 5549 5321 5583 5355
rect 14381 5321 14415 5355
rect 19901 5321 19935 5355
rect 20729 5321 20763 5355
rect 4997 5253 5031 5287
rect 10517 5253 10551 5287
rect 17785 5253 17819 5287
rect 18061 5253 18095 5287
rect 4629 5185 4663 5219
rect 4813 5185 4847 5219
rect 5457 5185 5491 5219
rect 8125 5185 8159 5219
rect 10701 5185 10735 5219
rect 14565 5185 14599 5219
rect 14749 5185 14783 5219
rect 15393 5185 15427 5219
rect 17877 5185 17911 5219
rect 20269 5185 20303 5219
rect 21097 5185 21131 5219
rect 23673 5185 23707 5219
rect 5641 5117 5675 5151
rect 8033 5117 8067 5151
rect 8493 5117 8527 5151
rect 8769 5117 8803 5151
rect 15301 5117 15335 5151
rect 15761 5117 15795 5151
rect 17417 5117 17451 5151
rect 17601 5117 17635 5151
rect 20361 5117 20395 5151
rect 20453 5117 20487 5151
rect 21189 5117 21223 5151
rect 21281 5117 21315 5151
rect 8953 5049 8987 5083
rect 10333 5049 10367 5083
rect 18245 5049 18279 5083
rect 23489 5049 23523 5083
rect 8585 4981 8619 5015
rect 5549 4777 5583 4811
rect 10885 4777 10919 4811
rect 11345 4777 11379 4811
rect 14933 4777 14967 4811
rect 20499 4777 20533 4811
rect 20867 4777 20901 4811
rect 7941 4709 7975 4743
rect 15301 4709 15335 4743
rect 4905 4641 4939 4675
rect 5825 4641 5859 4675
rect 7849 4641 7883 4675
rect 10609 4641 10643 4675
rect 10977 4641 11011 4675
rect 22477 4641 22511 4675
rect 5917 4573 5951 4607
rect 7665 4573 7699 4607
rect 8125 4573 8159 4607
rect 10517 4573 10551 4607
rect 11161 4573 11195 4607
rect 15117 4573 15151 4607
rect 20602 4573 20636 4607
rect 20796 4573 20830 4607
rect 23673 4573 23707 4607
rect 5089 4505 5123 4539
rect 7481 4505 7515 4539
rect 4997 4437 5031 4471
rect 5457 4437 5491 4471
rect 8309 4437 8343 4471
rect 4537 4233 4571 4267
rect 5273 4233 5307 4267
rect 7021 4233 7055 4267
rect 8125 4233 8159 4267
rect 10057 4165 10091 4199
rect 10241 4165 10275 4199
rect 3709 4097 3743 4131
rect 4813 4097 4847 4131
rect 5457 4097 5491 4131
rect 7297 4097 7331 4131
rect 10701 4097 10735 4131
rect 14381 4097 14415 4131
rect 15209 4097 15243 4131
rect 16037 4097 16071 4131
rect 17601 4097 17635 4131
rect 18429 4097 18463 4131
rect 3893 4029 3927 4063
rect 4353 4029 4387 4063
rect 4721 4029 4755 4063
rect 5181 4029 5215 4063
rect 5641 4029 5675 4063
rect 6653 4029 6687 4063
rect 6837 4029 6871 4063
rect 7389 4029 7423 4063
rect 7665 4029 7699 4063
rect 7849 4029 7883 4063
rect 8033 4029 8067 4063
rect 9873 4029 9907 4063
rect 10793 4029 10827 4063
rect 10885 4029 10919 4063
rect 14473 4029 14507 4063
rect 14749 4029 14783 4063
rect 15025 4029 15059 4063
rect 15117 4029 15151 4063
rect 15853 4029 15887 4063
rect 17693 4029 17727 4063
rect 17877 4029 17911 4063
rect 18061 4029 18095 4063
rect 18337 4029 18371 4063
rect 4077 3961 4111 3995
rect 4169 3961 4203 3995
rect 8493 3961 8527 3995
rect 10333 3961 10367 3995
rect 15577 3961 15611 3995
rect 15669 3961 15703 3995
rect 17233 3961 17267 3995
rect 4997 3689 5031 3723
rect 7941 3689 7975 3723
rect 10609 3689 10643 3723
rect 10701 3689 10735 3723
rect 14749 3689 14783 3723
rect 15209 3689 15243 3723
rect 16865 3689 16899 3723
rect 17785 3689 17819 3723
rect 18337 3689 18371 3723
rect 23489 3689 23523 3723
rect 11069 3621 11103 3655
rect 11529 3621 11563 3655
rect 17233 3621 17267 3655
rect 17325 3621 17359 3655
rect 10057 3553 10091 3587
rect 10885 3553 10919 3587
rect 12081 3553 12115 3587
rect 14381 3553 14415 3587
rect 17693 3553 17727 3587
rect 18981 3553 19015 3587
rect 4629 3485 4663 3519
rect 7573 3485 7607 3519
rect 7757 3485 7791 3519
rect 12474 3485 12508 3519
rect 14565 3485 14599 3519
rect 15025 3485 15059 3519
rect 17049 3485 17083 3519
rect 17509 3485 17543 3519
rect 17969 3485 18003 3519
rect 23673 3485 23707 3519
rect 4813 3417 4847 3451
rect 10241 3417 10275 3451
rect 14841 3417 14875 3451
rect 18153 3417 18187 3451
rect 18705 3417 18739 3451
rect 10149 3349 10183 3383
rect 11897 3349 11931 3383
rect 11989 3349 12023 3383
rect 12403 3349 12437 3383
rect 18797 3349 18831 3383
rect 4813 3145 4847 3179
rect 6653 3145 6687 3179
rect 7021 3145 7055 3179
rect 7481 3145 7515 3179
rect 10287 3145 10321 3179
rect 14657 3145 14691 3179
rect 15485 3145 15519 3179
rect 17693 3145 17727 3179
rect 18843 3145 18877 3179
rect 23489 3145 23523 3179
rect 5181 3077 5215 3111
rect 7849 3077 7883 3111
rect 18061 3077 18095 3111
rect 4572 3009 4606 3043
rect 5273 3009 5307 3043
rect 5687 3009 5721 3043
rect 5790 3009 5824 3043
rect 7941 3009 7975 3043
rect 8355 3009 8389 3043
rect 8458 3009 8492 3043
rect 10184 3009 10218 3043
rect 15025 3009 15059 3043
rect 15853 3009 15887 3043
rect 18153 3009 18187 3043
rect 18567 3009 18601 3043
rect 18670 3009 18704 3043
rect 18946 3009 18980 3043
rect 23673 3009 23707 3043
rect 5365 2941 5399 2975
rect 7113 2941 7147 2975
rect 7205 2941 7239 2975
rect 8033 2941 8067 2975
rect 15117 2941 15151 2975
rect 15301 2941 15335 2975
rect 15945 2941 15979 2975
rect 16129 2941 16163 2975
rect 18337 2941 18371 2975
rect 4675 2805 4709 2839
rect 4169 2601 4203 2635
rect 4537 2601 4571 2635
rect 4629 2601 4663 2635
rect 6101 2601 6135 2635
rect 7435 2601 7469 2635
rect 10609 2601 10643 2635
rect 11253 2601 11287 2635
rect 11897 2601 11931 2635
rect 12541 2601 12575 2635
rect 13185 2601 13219 2635
rect 14289 2601 14323 2635
rect 14979 2601 15013 2635
rect 15347 2601 15381 2635
rect 18797 2601 18831 2635
rect 19441 2601 19475 2635
rect 21373 2601 21407 2635
rect 5641 2533 5675 2567
rect 7297 2533 7331 2567
rect 15485 2533 15519 2567
rect 17509 2533 17543 2567
rect 5089 2465 5123 2499
rect 5273 2465 5307 2499
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4353 2397 4387 2431
rect 4997 2397 5031 2431
rect 5457 2397 5491 2431
rect 5917 2397 5951 2431
rect 6745 2397 6779 2431
rect 7113 2397 7147 2431
rect 7506 2397 7540 2431
rect 8033 2397 8067 2431
rect 8677 2397 8711 2431
rect 9321 2397 9355 2431
rect 9965 2397 9999 2431
rect 10425 2397 10459 2431
rect 11069 2397 11103 2431
rect 11713 2397 11747 2431
rect 12357 2397 12391 2431
rect 13001 2397 13035 2431
rect 13829 2397 13863 2431
rect 14473 2397 14507 2431
rect 15050 2397 15084 2431
rect 15276 2397 15310 2431
rect 15669 2397 15703 2431
rect 15945 2397 15979 2431
rect 16405 2397 16439 2431
rect 17049 2397 17083 2431
rect 17693 2397 17727 2431
rect 18337 2397 18371 2431
rect 18981 2397 19015 2431
rect 19625 2397 19659 2431
rect 20269 2397 20303 2431
rect 20913 2397 20947 2431
rect 21557 2397 21591 2431
rect 3525 2261 3559 2295
rect 6561 2261 6595 2295
rect 7849 2261 7883 2295
rect 8493 2261 8527 2295
rect 9137 2261 9171 2295
rect 9781 2261 9815 2295
rect 13645 2261 13679 2295
rect 15761 2261 15795 2295
rect 16221 2261 16255 2295
rect 16865 2261 16899 2295
rect 18153 2261 18187 2295
rect 20085 2261 20119 2295
rect 20729 2261 20763 2295
<< metal1 >>
rect 1104 25050 24012 25072
rect 1104 24998 4473 25050
rect 4525 24998 4537 25050
rect 4589 24998 4601 25050
rect 4653 24998 4665 25050
rect 4717 24998 4729 25050
rect 4781 24998 10200 25050
rect 10252 24998 10264 25050
rect 10316 24998 10328 25050
rect 10380 24998 10392 25050
rect 10444 24998 10456 25050
rect 10508 24998 15927 25050
rect 15979 24998 15991 25050
rect 16043 24998 16055 25050
rect 16107 24998 16119 25050
rect 16171 24998 16183 25050
rect 16235 24998 21654 25050
rect 21706 24998 21718 25050
rect 21770 24998 21782 25050
rect 21834 24998 21846 25050
rect 21898 24998 21910 25050
rect 21962 24998 24012 25050
rect 1104 24976 24012 24998
rect 5810 24760 5816 24812
rect 5868 24800 5874 24812
rect 5905 24803 5963 24809
rect 5905 24800 5917 24803
rect 5868 24772 5917 24800
rect 5868 24760 5874 24772
rect 5905 24769 5917 24772
rect 5951 24769 5963 24803
rect 5905 24763 5963 24769
rect 6454 24760 6460 24812
rect 6512 24800 6518 24812
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 6512 24772 6561 24800
rect 6512 24760 6518 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 7098 24760 7104 24812
rect 7156 24800 7162 24812
rect 7193 24803 7251 24809
rect 7193 24800 7205 24803
rect 7156 24772 7205 24800
rect 7156 24760 7162 24772
rect 7193 24769 7205 24772
rect 7239 24769 7251 24803
rect 7193 24763 7251 24769
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 7837 24803 7895 24809
rect 7837 24800 7849 24803
rect 7800 24772 7849 24800
rect 7800 24760 7806 24772
rect 7837 24769 7849 24772
rect 7883 24769 7895 24803
rect 7837 24763 7895 24769
rect 8662 24760 8668 24812
rect 8720 24760 8726 24812
rect 9122 24760 9128 24812
rect 9180 24800 9186 24812
rect 9309 24803 9367 24809
rect 9309 24800 9321 24803
rect 9180 24772 9321 24800
rect 9180 24760 9186 24772
rect 9309 24769 9321 24772
rect 9355 24769 9367 24803
rect 9309 24763 9367 24769
rect 9858 24760 9864 24812
rect 9916 24800 9922 24812
rect 9953 24803 10011 24809
rect 9953 24800 9965 24803
rect 9916 24772 9965 24800
rect 9916 24760 9922 24772
rect 9953 24769 9965 24772
rect 9999 24769 10011 24803
rect 9953 24763 10011 24769
rect 10042 24760 10048 24812
rect 10100 24800 10106 24812
rect 10597 24803 10655 24809
rect 10597 24800 10609 24803
rect 10100 24772 10609 24800
rect 10100 24760 10106 24772
rect 10597 24769 10609 24772
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 11054 24760 11060 24812
rect 11112 24800 11118 24812
rect 11241 24803 11299 24809
rect 11241 24800 11253 24803
rect 11112 24772 11253 24800
rect 11112 24760 11118 24772
rect 11241 24769 11253 24772
rect 11287 24769 11299 24803
rect 11241 24763 11299 24769
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 11664 24772 11713 24800
rect 11664 24760 11670 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 12250 24760 12256 24812
rect 12308 24800 12314 24812
rect 12345 24803 12403 24809
rect 12345 24800 12357 24803
rect 12308 24772 12357 24800
rect 12308 24760 12314 24772
rect 12345 24769 12357 24772
rect 12391 24769 12403 24803
rect 12345 24763 12403 24769
rect 12894 24760 12900 24812
rect 12952 24800 12958 24812
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12952 24772 13001 24800
rect 12952 24760 12958 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13538 24760 13544 24812
rect 13596 24800 13602 24812
rect 13817 24803 13875 24809
rect 13817 24800 13829 24803
rect 13596 24772 13829 24800
rect 13596 24760 13602 24772
rect 13817 24769 13829 24772
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 14458 24760 14464 24812
rect 14516 24760 14522 24812
rect 14826 24760 14832 24812
rect 14884 24800 14890 24812
rect 15105 24803 15163 24809
rect 15105 24800 15117 24803
rect 14884 24772 15117 24800
rect 14884 24760 14890 24772
rect 15105 24769 15117 24772
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 15746 24760 15752 24812
rect 15804 24760 15810 24812
rect 16390 24760 16396 24812
rect 16448 24760 16454 24812
rect 16758 24760 16764 24812
rect 16816 24800 16822 24812
rect 17037 24803 17095 24809
rect 17037 24800 17049 24803
rect 16816 24772 17049 24800
rect 16816 24760 16822 24772
rect 17037 24769 17049 24772
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 17497 24803 17555 24809
rect 17497 24800 17509 24803
rect 17460 24772 17509 24800
rect 17460 24760 17466 24772
rect 17497 24769 17509 24772
rect 17543 24769 17555 24803
rect 17497 24763 17555 24769
rect 18046 24760 18052 24812
rect 18104 24800 18110 24812
rect 18141 24803 18199 24809
rect 18141 24800 18153 24803
rect 18104 24772 18153 24800
rect 18104 24760 18110 24772
rect 18141 24769 18153 24772
rect 18187 24769 18199 24803
rect 18141 24763 18199 24769
rect 20622 24760 20628 24812
rect 20680 24800 20686 24812
rect 20717 24803 20775 24809
rect 20717 24800 20729 24803
rect 20680 24772 20729 24800
rect 20680 24760 20686 24772
rect 20717 24769 20729 24772
rect 20763 24769 20775 24803
rect 20717 24763 20775 24769
rect 23658 24760 23664 24812
rect 23716 24760 23722 24812
rect 22738 24692 22744 24744
rect 22796 24692 22802 24744
rect 8386 24624 8392 24676
rect 8444 24664 8450 24676
rect 8481 24667 8539 24673
rect 8481 24664 8493 24667
rect 8444 24636 8493 24664
rect 8444 24624 8450 24636
rect 8481 24633 8493 24636
rect 8527 24633 8539 24667
rect 8481 24627 8539 24633
rect 9030 24624 9036 24676
rect 9088 24664 9094 24676
rect 9125 24667 9183 24673
rect 9125 24664 9137 24667
rect 9088 24636 9137 24664
rect 9088 24624 9094 24636
rect 9125 24633 9137 24636
rect 9171 24633 9183 24667
rect 9125 24627 9183 24633
rect 9674 24624 9680 24676
rect 9732 24664 9738 24676
rect 9769 24667 9827 24673
rect 9769 24664 9781 24667
rect 9732 24636 9781 24664
rect 9732 24624 9738 24636
rect 9769 24633 9781 24636
rect 9815 24633 9827 24667
rect 9769 24627 9827 24633
rect 10413 24667 10471 24673
rect 10413 24633 10425 24667
rect 10459 24664 10471 24667
rect 10594 24664 10600 24676
rect 10459 24636 10600 24664
rect 10459 24633 10471 24636
rect 10413 24627 10471 24633
rect 10594 24624 10600 24636
rect 10652 24624 10658 24676
rect 10962 24624 10968 24676
rect 11020 24664 11026 24676
rect 11057 24667 11115 24673
rect 11057 24664 11069 24667
rect 11020 24636 11069 24664
rect 11020 24624 11026 24636
rect 11057 24633 11069 24636
rect 11103 24633 11115 24667
rect 11057 24627 11115 24633
rect 14182 24624 14188 24676
rect 14240 24664 14246 24676
rect 14277 24667 14335 24673
rect 14277 24664 14289 24667
rect 14240 24636 14289 24664
rect 14240 24624 14246 24636
rect 14277 24633 14289 24636
rect 14323 24633 14335 24667
rect 14277 24627 14335 24633
rect 15470 24624 15476 24676
rect 15528 24664 15534 24676
rect 15565 24667 15623 24673
rect 15565 24664 15577 24667
rect 15528 24636 15577 24664
rect 15528 24624 15534 24636
rect 15565 24633 15577 24636
rect 15611 24633 15623 24667
rect 15565 24627 15623 24633
rect 16209 24667 16267 24673
rect 16209 24633 16221 24667
rect 16255 24664 16267 24667
rect 16298 24664 16304 24676
rect 16255 24636 16304 24664
rect 16255 24633 16267 24636
rect 16209 24627 16267 24633
rect 16298 24624 16304 24636
rect 16356 24624 16362 24676
rect 6086 24556 6092 24608
rect 6144 24556 6150 24608
rect 6730 24556 6736 24608
rect 6788 24556 6794 24608
rect 7374 24556 7380 24608
rect 7432 24556 7438 24608
rect 8021 24599 8079 24605
rect 8021 24565 8033 24599
rect 8067 24596 8079 24599
rect 9306 24596 9312 24608
rect 8067 24568 9312 24596
rect 8067 24565 8079 24568
rect 8021 24559 8079 24565
rect 9306 24556 9312 24568
rect 9364 24556 9370 24608
rect 11882 24556 11888 24608
rect 11940 24556 11946 24608
rect 12526 24556 12532 24608
rect 12584 24556 12590 24608
rect 12802 24556 12808 24608
rect 12860 24596 12866 24608
rect 13173 24599 13231 24605
rect 13173 24596 13185 24599
rect 12860 24568 13185 24596
rect 12860 24556 12866 24568
rect 13173 24565 13185 24568
rect 13219 24565 13231 24599
rect 13173 24559 13231 24565
rect 13630 24556 13636 24608
rect 13688 24556 13694 24608
rect 14918 24556 14924 24608
rect 14976 24556 14982 24608
rect 16850 24556 16856 24608
rect 16908 24556 16914 24608
rect 17586 24556 17592 24608
rect 17644 24596 17650 24608
rect 17681 24599 17739 24605
rect 17681 24596 17693 24599
rect 17644 24568 17693 24596
rect 17644 24556 17650 24568
rect 17681 24565 17693 24568
rect 17727 24565 17739 24599
rect 17681 24559 17739 24565
rect 18322 24556 18328 24608
rect 18380 24556 18386 24608
rect 20898 24556 20904 24608
rect 20956 24556 20962 24608
rect 1104 24506 24012 24528
rect 1104 24454 3813 24506
rect 3865 24454 3877 24506
rect 3929 24454 3941 24506
rect 3993 24454 4005 24506
rect 4057 24454 4069 24506
rect 4121 24454 9540 24506
rect 9592 24454 9604 24506
rect 9656 24454 9668 24506
rect 9720 24454 9732 24506
rect 9784 24454 9796 24506
rect 9848 24454 15267 24506
rect 15319 24454 15331 24506
rect 15383 24454 15395 24506
rect 15447 24454 15459 24506
rect 15511 24454 15523 24506
rect 15575 24454 20994 24506
rect 21046 24454 21058 24506
rect 21110 24454 21122 24506
rect 21174 24454 21186 24506
rect 21238 24454 21250 24506
rect 21302 24454 24012 24506
rect 1104 24432 24012 24454
rect 23014 24216 23020 24268
rect 23072 24216 23078 24268
rect 7374 24148 7380 24200
rect 7432 24188 7438 24200
rect 9058 24191 9116 24197
rect 9058 24188 9070 24191
rect 7432 24160 9070 24188
rect 7432 24148 7438 24160
rect 9058 24157 9070 24160
rect 9104 24157 9116 24191
rect 9058 24151 9116 24157
rect 14804 24191 14862 24197
rect 14804 24157 14816 24191
rect 14850 24188 14862 24191
rect 16850 24188 16856 24200
rect 14850 24160 16856 24188
rect 14850 24157 14862 24160
rect 14804 24151 14862 24157
rect 16850 24148 16856 24160
rect 16908 24148 16914 24200
rect 23658 24148 23664 24200
rect 23716 24148 23722 24200
rect 8386 24012 8392 24064
rect 8444 24052 8450 24064
rect 8987 24055 9045 24061
rect 8987 24052 8999 24055
rect 8444 24024 8999 24052
rect 8444 24012 8450 24024
rect 8987 24021 8999 24024
rect 9033 24021 9045 24055
rect 8987 24015 9045 24021
rect 14875 24055 14933 24061
rect 14875 24021 14887 24055
rect 14921 24052 14933 24055
rect 15562 24052 15568 24064
rect 14921 24024 15568 24052
rect 14921 24021 14933 24024
rect 14875 24015 14933 24021
rect 15562 24012 15568 24024
rect 15620 24012 15626 24064
rect 1104 23962 24012 23984
rect 1104 23910 4473 23962
rect 4525 23910 4537 23962
rect 4589 23910 4601 23962
rect 4653 23910 4665 23962
rect 4717 23910 4729 23962
rect 4781 23910 10200 23962
rect 10252 23910 10264 23962
rect 10316 23910 10328 23962
rect 10380 23910 10392 23962
rect 10444 23910 10456 23962
rect 10508 23910 15927 23962
rect 15979 23910 15991 23962
rect 16043 23910 16055 23962
rect 16107 23910 16119 23962
rect 16171 23910 16183 23962
rect 16235 23910 21654 23962
rect 21706 23910 21718 23962
rect 21770 23910 21782 23962
rect 21834 23910 21846 23962
rect 21898 23910 21910 23962
rect 21962 23910 24012 23962
rect 1104 23888 24012 23910
rect 8386 23808 8392 23860
rect 8444 23808 8450 23860
rect 9306 23808 9312 23860
rect 9364 23808 9370 23860
rect 14645 23851 14703 23857
rect 14645 23817 14657 23851
rect 14691 23848 14703 23851
rect 14918 23848 14924 23860
rect 14691 23820 14924 23848
rect 14691 23817 14703 23820
rect 14645 23811 14703 23817
rect 14918 23808 14924 23820
rect 14976 23808 14982 23860
rect 15562 23808 15568 23860
rect 15620 23808 15626 23860
rect 17586 23808 17592 23860
rect 17644 23848 17650 23860
rect 17644 23820 18276 23848
rect 17644 23808 17650 23820
rect 7374 23740 7380 23792
rect 7432 23780 7438 23792
rect 8481 23783 8539 23789
rect 8481 23780 8493 23783
rect 7432 23752 8493 23780
rect 7432 23740 7438 23752
rect 8481 23749 8493 23752
rect 8527 23749 8539 23783
rect 9324 23780 9352 23808
rect 15473 23783 15531 23789
rect 9324 23752 9996 23780
rect 8481 23743 8539 23749
rect 9968 23721 9996 23752
rect 15473 23749 15485 23783
rect 15519 23780 15531 23783
rect 16850 23780 16856 23792
rect 15519 23752 16856 23780
rect 15519 23749 15531 23752
rect 15473 23743 15531 23749
rect 16850 23740 16856 23752
rect 16908 23740 16914 23792
rect 9401 23715 9459 23721
rect 9401 23681 9413 23715
rect 9447 23712 9459 23715
rect 9815 23715 9873 23721
rect 9815 23712 9827 23715
rect 9447 23684 9827 23712
rect 9447 23681 9459 23684
rect 9401 23675 9459 23681
rect 9815 23681 9827 23684
rect 9861 23681 9873 23715
rect 9815 23675 9873 23681
rect 9918 23715 9996 23721
rect 9918 23681 9930 23715
rect 9964 23684 9996 23715
rect 9964 23681 9976 23684
rect 9918 23675 9976 23681
rect 12342 23672 12348 23724
rect 12400 23712 12406 23724
rect 18248 23721 18276 23820
rect 17681 23715 17739 23721
rect 12400 23684 16574 23712
rect 12400 23672 12406 23684
rect 8294 23604 8300 23656
rect 8352 23644 8358 23656
rect 8352 23616 8708 23644
rect 8352 23604 8358 23616
rect 8680 23576 8708 23616
rect 8754 23604 8760 23656
rect 8812 23644 8818 23656
rect 9493 23647 9551 23653
rect 9493 23644 9505 23647
rect 8812 23616 9505 23644
rect 8812 23604 8818 23616
rect 9493 23613 9505 23616
rect 9539 23613 9551 23647
rect 9493 23607 9551 23613
rect 14734 23604 14740 23656
rect 14792 23604 14798 23656
rect 14936 23653 14964 23684
rect 14921 23647 14979 23653
rect 14921 23613 14933 23647
rect 14967 23613 14979 23647
rect 14921 23607 14979 23613
rect 15654 23604 15660 23656
rect 15712 23604 15718 23656
rect 16546 23644 16574 23684
rect 17681 23681 17693 23715
rect 17727 23712 17739 23715
rect 18095 23715 18153 23721
rect 18095 23712 18107 23715
rect 17727 23684 18107 23712
rect 17727 23681 17739 23684
rect 17681 23675 17739 23681
rect 18095 23681 18107 23684
rect 18141 23681 18153 23715
rect 18095 23675 18153 23681
rect 18198 23715 18276 23721
rect 18198 23681 18210 23715
rect 18244 23684 18276 23715
rect 18244 23681 18256 23684
rect 18198 23675 18256 23681
rect 18322 23672 18328 23724
rect 18380 23712 18386 23724
rect 18442 23715 18500 23721
rect 18442 23712 18454 23715
rect 18380 23684 18454 23712
rect 18380 23672 18386 23684
rect 18442 23681 18454 23684
rect 18488 23681 18500 23715
rect 18442 23675 18500 23681
rect 23382 23672 23388 23724
rect 23440 23712 23446 23724
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 23440 23684 23673 23712
rect 23440 23672 23446 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 17865 23647 17923 23653
rect 17865 23644 17877 23647
rect 16546 23616 17877 23644
rect 17865 23613 17877 23616
rect 17911 23644 17923 23647
rect 20622 23644 20628 23656
rect 17911 23616 20628 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 20622 23604 20628 23616
rect 20680 23604 20686 23656
rect 12342 23576 12348 23588
rect 8680 23548 12348 23576
rect 12342 23536 12348 23548
rect 12400 23536 12406 23588
rect 8846 23468 8852 23520
rect 8904 23468 8910 23520
rect 8941 23511 8999 23517
rect 8941 23477 8953 23511
rect 8987 23508 8999 23511
rect 9030 23508 9036 23520
rect 8987 23480 9036 23508
rect 8987 23477 8999 23480
rect 8941 23471 8999 23477
rect 9030 23468 9036 23480
rect 9088 23468 9094 23520
rect 14274 23468 14280 23520
rect 14332 23468 14338 23520
rect 15010 23468 15016 23520
rect 15068 23508 15074 23520
rect 15105 23511 15163 23517
rect 15105 23508 15117 23511
rect 15068 23480 15117 23508
rect 15068 23468 15074 23480
rect 15105 23477 15117 23480
rect 15151 23477 15163 23511
rect 15105 23471 15163 23477
rect 17034 23468 17040 23520
rect 17092 23508 17098 23520
rect 17221 23511 17279 23517
rect 17221 23508 17233 23511
rect 17092 23480 17233 23508
rect 17092 23468 17098 23480
rect 17221 23477 17233 23480
rect 17267 23477 17279 23511
rect 17221 23471 17279 23477
rect 18046 23468 18052 23520
rect 18104 23508 18110 23520
rect 18371 23511 18429 23517
rect 18371 23508 18383 23511
rect 18104 23480 18383 23508
rect 18104 23468 18110 23480
rect 18371 23477 18383 23480
rect 18417 23477 18429 23511
rect 18371 23471 18429 23477
rect 23477 23511 23535 23517
rect 23477 23477 23489 23511
rect 23523 23508 23535 23511
rect 23842 23508 23848 23520
rect 23523 23480 23848 23508
rect 23523 23477 23535 23480
rect 23477 23471 23535 23477
rect 23842 23468 23848 23480
rect 23900 23468 23906 23520
rect 1104 23418 24012 23440
rect 1104 23366 3813 23418
rect 3865 23366 3877 23418
rect 3929 23366 3941 23418
rect 3993 23366 4005 23418
rect 4057 23366 4069 23418
rect 4121 23366 9540 23418
rect 9592 23366 9604 23418
rect 9656 23366 9668 23418
rect 9720 23366 9732 23418
rect 9784 23366 9796 23418
rect 9848 23366 15267 23418
rect 15319 23366 15331 23418
rect 15383 23366 15395 23418
rect 15447 23366 15459 23418
rect 15511 23366 15523 23418
rect 15575 23366 20994 23418
rect 21046 23366 21058 23418
rect 21110 23366 21122 23418
rect 21174 23366 21186 23418
rect 21238 23366 21250 23418
rect 21302 23366 24012 23418
rect 1104 23344 24012 23366
rect 14734 23313 14740 23316
rect 14691 23307 14740 23313
rect 14691 23273 14703 23307
rect 14737 23273 14740 23307
rect 14691 23267 14740 23273
rect 14734 23264 14740 23267
rect 14792 23264 14798 23316
rect 6822 23128 6828 23180
rect 6880 23168 6886 23180
rect 6917 23171 6975 23177
rect 6917 23168 6929 23171
rect 6880 23140 6929 23168
rect 6880 23128 6886 23140
rect 6917 23137 6929 23140
rect 6963 23137 6975 23171
rect 6917 23131 6975 23137
rect 15654 23128 15660 23180
rect 15712 23168 15718 23180
rect 17957 23171 18015 23177
rect 17957 23168 17969 23171
rect 15712 23140 17969 23168
rect 15712 23128 15718 23140
rect 17957 23137 17969 23140
rect 18003 23168 18015 23171
rect 22738 23168 22744 23180
rect 18003 23140 22744 23168
rect 18003 23137 18015 23140
rect 17957 23131 18015 23137
rect 22738 23128 22744 23140
rect 22796 23128 22802 23180
rect 6086 23060 6092 23112
rect 6144 23100 6150 23112
rect 6733 23103 6791 23109
rect 6733 23100 6745 23103
rect 6144 23072 6745 23100
rect 6144 23060 6150 23072
rect 6733 23069 6745 23072
rect 6779 23100 6791 23103
rect 7310 23103 7368 23109
rect 7310 23100 7322 23103
rect 6779 23072 7322 23100
rect 6779 23069 6791 23072
rect 6733 23063 6791 23069
rect 7310 23069 7322 23072
rect 7356 23069 7368 23103
rect 7310 23063 7368 23069
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8904 23072 8953 23100
rect 8904 23060 8910 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 9088 23072 9137 23100
rect 9088 23060 9094 23072
rect 9125 23069 9137 23072
rect 9171 23069 9183 23103
rect 9125 23063 9183 23069
rect 14794 23103 14852 23109
rect 14794 23069 14806 23103
rect 14840 23100 14852 23103
rect 14918 23100 14924 23112
rect 14840 23072 14924 23100
rect 14840 23069 14852 23072
rect 14794 23063 14852 23069
rect 14918 23060 14924 23072
rect 14976 23060 14982 23112
rect 17865 23103 17923 23109
rect 17865 23069 17877 23103
rect 17911 23100 17923 23103
rect 18046 23100 18052 23112
rect 17911 23072 18052 23100
rect 17911 23069 17923 23072
rect 17865 23063 17923 23069
rect 18046 23060 18052 23072
rect 18104 23060 18110 23112
rect 17773 23035 17831 23041
rect 17773 23001 17785 23035
rect 17819 23032 17831 23035
rect 18322 23032 18328 23044
rect 17819 23004 18328 23032
rect 17819 23001 17831 23004
rect 17773 22995 17831 23001
rect 18322 22992 18328 23004
rect 18380 22992 18386 23044
rect 6362 22924 6368 22976
rect 6420 22924 6426 22976
rect 6825 22967 6883 22973
rect 6825 22933 6837 22967
rect 6871 22964 6883 22967
rect 7239 22967 7297 22973
rect 7239 22964 7251 22967
rect 6871 22936 7251 22964
rect 6871 22933 6883 22936
rect 6825 22927 6883 22933
rect 7239 22933 7251 22936
rect 7285 22933 7297 22967
rect 7239 22927 7297 22933
rect 9309 22967 9367 22973
rect 9309 22933 9321 22967
rect 9355 22964 9367 22967
rect 9490 22964 9496 22976
rect 9355 22936 9496 22964
rect 9355 22933 9367 22936
rect 9309 22927 9367 22933
rect 9490 22924 9496 22936
rect 9548 22924 9554 22976
rect 17402 22924 17408 22976
rect 17460 22924 17466 22976
rect 1104 22874 24012 22896
rect 1104 22822 4473 22874
rect 4525 22822 4537 22874
rect 4589 22822 4601 22874
rect 4653 22822 4665 22874
rect 4717 22822 4729 22874
rect 4781 22822 10200 22874
rect 10252 22822 10264 22874
rect 10316 22822 10328 22874
rect 10380 22822 10392 22874
rect 10444 22822 10456 22874
rect 10508 22822 15927 22874
rect 15979 22822 15991 22874
rect 16043 22822 16055 22874
rect 16107 22822 16119 22874
rect 16171 22822 16183 22874
rect 16235 22822 21654 22874
rect 21706 22822 21718 22874
rect 21770 22822 21782 22874
rect 21834 22822 21846 22874
rect 21898 22822 21910 22874
rect 21962 22822 24012 22874
rect 1104 22800 24012 22822
rect 6917 22763 6975 22769
rect 6917 22729 6929 22763
rect 6963 22760 6975 22763
rect 7331 22763 7389 22769
rect 7331 22760 7343 22763
rect 6963 22732 7343 22760
rect 6963 22729 6975 22732
rect 6917 22723 6975 22729
rect 7331 22729 7343 22732
rect 7377 22729 7389 22763
rect 7331 22723 7389 22729
rect 9490 22720 9496 22772
rect 9548 22720 9554 22772
rect 11882 22720 11888 22772
rect 11940 22760 11946 22772
rect 12069 22763 12127 22769
rect 12069 22760 12081 22763
rect 11940 22732 12081 22760
rect 11940 22720 11946 22732
rect 12069 22729 12081 22732
rect 12115 22729 12127 22763
rect 12069 22723 12127 22729
rect 20441 22763 20499 22769
rect 20441 22729 20453 22763
rect 20487 22760 20499 22763
rect 20898 22760 20904 22772
rect 20487 22732 20904 22760
rect 20487 22729 20499 22732
rect 20441 22723 20499 22729
rect 12084 22692 12112 22723
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 14921 22695 14979 22701
rect 14921 22692 14933 22695
rect 6840 22664 7144 22692
rect 12084 22664 12756 22692
rect 6730 22584 6736 22636
rect 6788 22624 6794 22636
rect 6840 22633 6868 22664
rect 6825 22627 6883 22633
rect 6825 22624 6837 22627
rect 6788 22596 6837 22624
rect 6788 22584 6794 22596
rect 6825 22593 6837 22596
rect 6871 22593 6883 22627
rect 7116 22624 7144 22664
rect 7402 22627 7460 22633
rect 7402 22624 7414 22627
rect 7116 22596 7414 22624
rect 6825 22587 6883 22593
rect 7402 22593 7414 22596
rect 7448 22593 7460 22627
rect 7402 22587 7460 22593
rect 8573 22627 8631 22633
rect 8573 22593 8585 22627
rect 8619 22624 8631 22627
rect 8846 22624 8852 22636
rect 8619 22596 8852 22624
rect 8619 22593 8631 22596
rect 8573 22587 8631 22593
rect 8846 22584 8852 22596
rect 8904 22584 8910 22636
rect 9398 22584 9404 22636
rect 9456 22584 9462 22636
rect 12728 22633 12756 22664
rect 14476 22664 14933 22692
rect 14476 22633 14504 22664
rect 14921 22661 14933 22664
rect 14967 22692 14979 22695
rect 15010 22692 15016 22704
rect 14967 22664 15016 22692
rect 14967 22661 14979 22664
rect 14921 22655 14979 22661
rect 15010 22652 15016 22664
rect 15068 22652 15074 22704
rect 20916 22692 20944 22720
rect 20916 22664 21128 22692
rect 10045 22627 10103 22633
rect 10045 22624 10057 22627
rect 9508 22596 10057 22624
rect 5534 22516 5540 22568
rect 5592 22556 5598 22568
rect 7101 22559 7159 22565
rect 7101 22556 7113 22559
rect 5592 22528 7113 22556
rect 5592 22516 5598 22528
rect 7101 22525 7113 22528
rect 7147 22556 7159 22559
rect 8294 22556 8300 22568
rect 7147 22528 8300 22556
rect 7147 22525 7159 22528
rect 7101 22519 7159 22525
rect 8294 22516 8300 22528
rect 8352 22516 8358 22568
rect 8665 22559 8723 22565
rect 8665 22525 8677 22559
rect 8711 22556 8723 22559
rect 9030 22556 9036 22568
rect 8711 22528 9036 22556
rect 8711 22525 8723 22528
rect 8665 22519 8723 22525
rect 9030 22516 9036 22528
rect 9088 22556 9094 22568
rect 9214 22556 9220 22568
rect 9088 22528 9220 22556
rect 9088 22516 9094 22528
rect 9214 22516 9220 22528
rect 9272 22556 9278 22568
rect 9508 22556 9536 22596
rect 10045 22593 10057 22596
rect 10091 22593 10103 22627
rect 10045 22587 10103 22593
rect 12161 22627 12219 22633
rect 12161 22593 12173 22627
rect 12207 22624 12219 22627
rect 12575 22627 12633 22633
rect 12575 22624 12587 22627
rect 12207 22596 12587 22624
rect 12207 22593 12219 22596
rect 12161 22587 12219 22593
rect 12575 22593 12587 22596
rect 12621 22593 12633 22627
rect 12575 22587 12633 22593
rect 12678 22627 12756 22633
rect 12678 22593 12690 22627
rect 12724 22596 12756 22627
rect 14461 22627 14519 22633
rect 12724 22593 12736 22596
rect 12678 22587 12736 22593
rect 14461 22593 14473 22627
rect 14507 22593 14519 22627
rect 14461 22587 14519 22593
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 17221 22627 17279 22633
rect 17221 22593 17233 22627
rect 17267 22624 17279 22627
rect 17402 22624 17408 22636
rect 17267 22596 17408 22624
rect 17267 22593 17279 22596
rect 17221 22587 17279 22593
rect 9272 22528 9536 22556
rect 9272 22516 9278 22528
rect 9582 22516 9588 22568
rect 9640 22516 9646 22568
rect 12342 22516 12348 22568
rect 12400 22516 12406 22568
rect 14274 22516 14280 22568
rect 14332 22556 14338 22568
rect 14918 22556 14924 22568
rect 14332 22528 14924 22556
rect 14332 22516 14338 22528
rect 14918 22516 14924 22528
rect 14976 22556 14982 22568
rect 15120 22556 15148 22587
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 21100 22633 21128 22664
rect 20533 22627 20591 22633
rect 20533 22593 20545 22627
rect 20579 22624 20591 22627
rect 20947 22627 21005 22633
rect 20947 22624 20959 22627
rect 20579 22596 20959 22624
rect 20579 22593 20591 22596
rect 20533 22587 20591 22593
rect 20947 22593 20959 22596
rect 20993 22593 21005 22627
rect 20947 22587 21005 22593
rect 21050 22627 21128 22633
rect 21050 22593 21062 22627
rect 21096 22596 21128 22627
rect 21096 22593 21108 22596
rect 21050 22587 21108 22593
rect 23658 22584 23664 22636
rect 23716 22584 23722 22636
rect 14976 22528 15148 22556
rect 14976 22516 14982 22528
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 17034 22556 17040 22568
rect 16816 22528 17040 22556
rect 16816 22516 16822 22528
rect 17034 22516 17040 22528
rect 17092 22516 17098 22568
rect 20622 22516 20628 22568
rect 20680 22556 20686 22568
rect 23014 22556 23020 22568
rect 20680 22528 23020 22556
rect 20680 22516 20686 22528
rect 23014 22516 23020 22528
rect 23072 22516 23078 22568
rect 8846 22448 8852 22500
rect 8904 22488 8910 22500
rect 9861 22491 9919 22497
rect 9861 22488 9873 22491
rect 8904 22460 9873 22488
rect 8904 22448 8910 22460
rect 9861 22457 9873 22460
rect 9907 22457 9919 22491
rect 9861 22451 9919 22457
rect 16666 22448 16672 22500
rect 16724 22488 16730 22500
rect 17494 22488 17500 22500
rect 16724 22460 17500 22488
rect 16724 22448 16730 22460
rect 17494 22448 17500 22460
rect 17552 22448 17558 22500
rect 6454 22380 6460 22432
rect 6512 22380 6518 22432
rect 8938 22380 8944 22432
rect 8996 22380 9002 22432
rect 9030 22380 9036 22432
rect 9088 22380 9094 22432
rect 9306 22380 9312 22432
rect 9364 22420 9370 22432
rect 9582 22420 9588 22432
rect 9364 22392 9588 22420
rect 9364 22380 9370 22392
rect 9582 22380 9588 22392
rect 9640 22380 9646 22432
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 10229 22423 10287 22429
rect 10229 22420 10241 22423
rect 10008 22392 10241 22420
rect 10008 22380 10014 22392
rect 10229 22389 10241 22392
rect 10275 22389 10287 22423
rect 10229 22383 10287 22389
rect 11701 22423 11759 22429
rect 11701 22389 11713 22423
rect 11747 22420 11759 22423
rect 11974 22420 11980 22432
rect 11747 22392 11980 22420
rect 11747 22389 11759 22392
rect 11701 22383 11759 22389
rect 11974 22380 11980 22392
rect 12032 22380 12038 22432
rect 14642 22380 14648 22432
rect 14700 22380 14706 22432
rect 14734 22380 14740 22432
rect 14792 22380 14798 22432
rect 17218 22380 17224 22432
rect 17276 22420 17282 22432
rect 17405 22423 17463 22429
rect 17405 22420 17417 22423
rect 17276 22392 17417 22420
rect 17276 22380 17282 22392
rect 17405 22389 17417 22392
rect 17451 22389 17463 22423
rect 17405 22383 17463 22389
rect 20073 22423 20131 22429
rect 20073 22389 20085 22423
rect 20119 22420 20131 22423
rect 20898 22420 20904 22432
rect 20119 22392 20904 22420
rect 20119 22389 20131 22392
rect 20073 22383 20131 22389
rect 20898 22380 20904 22392
rect 20956 22380 20962 22432
rect 23106 22380 23112 22432
rect 23164 22420 23170 22432
rect 23477 22423 23535 22429
rect 23477 22420 23489 22423
rect 23164 22392 23489 22420
rect 23164 22380 23170 22392
rect 23477 22389 23489 22392
rect 23523 22389 23535 22423
rect 23477 22383 23535 22389
rect 1104 22330 24012 22352
rect 1104 22278 3813 22330
rect 3865 22278 3877 22330
rect 3929 22278 3941 22330
rect 3993 22278 4005 22330
rect 4057 22278 4069 22330
rect 4121 22278 9540 22330
rect 9592 22278 9604 22330
rect 9656 22278 9668 22330
rect 9720 22278 9732 22330
rect 9784 22278 9796 22330
rect 9848 22278 15267 22330
rect 15319 22278 15331 22330
rect 15383 22278 15395 22330
rect 15447 22278 15459 22330
rect 15511 22278 15523 22330
rect 15575 22278 20994 22330
rect 21046 22278 21058 22330
rect 21110 22278 21122 22330
rect 21174 22278 21186 22330
rect 21238 22278 21250 22330
rect 21302 22278 24012 22330
rect 1104 22256 24012 22278
rect 5902 22176 5908 22228
rect 5960 22216 5966 22228
rect 6822 22216 6828 22228
rect 5960 22188 6828 22216
rect 5960 22176 5966 22188
rect 6822 22176 6828 22188
rect 6880 22216 6886 22228
rect 8754 22216 8760 22228
rect 6880 22188 8760 22216
rect 6880 22176 6886 22188
rect 8754 22176 8760 22188
rect 8812 22216 8818 22228
rect 9309 22219 9367 22225
rect 8812 22188 9260 22216
rect 8812 22176 8818 22188
rect 8846 22108 8852 22160
rect 8904 22148 8910 22160
rect 8941 22151 8999 22157
rect 8941 22148 8953 22151
rect 8904 22120 8953 22148
rect 8904 22108 8910 22120
rect 8941 22117 8953 22120
rect 8987 22117 8999 22151
rect 9232 22148 9260 22188
rect 9309 22185 9321 22219
rect 9355 22216 9367 22219
rect 9398 22216 9404 22228
rect 9355 22188 9404 22216
rect 9355 22185 9367 22188
rect 9309 22179 9367 22185
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 15654 22216 15660 22228
rect 12636 22188 15660 22216
rect 12636 22148 12664 22188
rect 15654 22176 15660 22188
rect 15712 22176 15718 22228
rect 17402 22176 17408 22228
rect 17460 22176 17466 22228
rect 9232 22120 12664 22148
rect 8941 22111 8999 22117
rect 9125 22083 9183 22089
rect 9125 22049 9137 22083
rect 9171 22080 9183 22083
rect 9214 22080 9220 22092
rect 9171 22052 9220 22080
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 9214 22040 9220 22052
rect 9272 22040 9278 22092
rect 12636 22089 12664 22120
rect 14844 22120 16528 22148
rect 14844 22089 14872 22120
rect 12621 22083 12679 22089
rect 12621 22080 12633 22083
rect 12599 22052 12633 22080
rect 12621 22049 12633 22052
rect 12667 22049 12679 22083
rect 12621 22043 12679 22049
rect 14829 22083 14887 22089
rect 14829 22049 14841 22083
rect 14875 22080 14887 22083
rect 14875 22052 14909 22080
rect 14875 22049 14887 22052
rect 14829 22043 14887 22049
rect 15010 22040 15016 22092
rect 15068 22040 15074 22092
rect 15102 22040 15108 22092
rect 15160 22080 15166 22092
rect 15289 22083 15347 22089
rect 15289 22080 15301 22083
rect 15160 22052 15301 22080
rect 15160 22040 15166 22052
rect 15289 22049 15301 22052
rect 15335 22049 15347 22083
rect 16500 22080 16528 22120
rect 16574 22108 16580 22160
rect 16632 22148 16638 22160
rect 17420 22148 17448 22176
rect 16632 22120 17816 22148
rect 16632 22108 16638 22120
rect 16666 22080 16672 22092
rect 16500 22052 16672 22080
rect 15289 22043 15347 22049
rect 16666 22040 16672 22052
rect 16724 22040 16730 22092
rect 17494 22040 17500 22092
rect 17552 22040 17558 22092
rect 17586 22040 17592 22092
rect 17644 22080 17650 22092
rect 17681 22083 17739 22089
rect 17681 22080 17693 22083
rect 17644 22052 17693 22080
rect 17644 22040 17650 22052
rect 17681 22049 17693 22052
rect 17727 22049 17739 22083
rect 17788 22080 17816 22120
rect 17957 22083 18015 22089
rect 17957 22080 17969 22083
rect 17788 22052 17969 22080
rect 17681 22043 17739 22049
rect 17957 22049 17969 22052
rect 18003 22049 18015 22083
rect 17957 22043 18015 22049
rect 6362 21972 6368 22024
rect 6420 22012 6426 22024
rect 12437 22015 12495 22021
rect 6420 21984 6684 22012
rect 6420 21972 6426 21984
rect 6656 21956 6684 21984
rect 12437 21981 12449 22015
rect 12483 22012 12495 22015
rect 12526 22012 12532 22024
rect 12483 21984 12532 22012
rect 12483 21981 12495 21984
rect 12437 21975 12495 21981
rect 12526 21972 12532 21984
rect 12584 22012 12590 22024
rect 13014 22015 13072 22021
rect 13014 22012 13026 22015
rect 12584 21984 13026 22012
rect 12584 21972 12590 21984
rect 13014 21981 13026 21984
rect 13060 21981 13072 22015
rect 13014 21975 13072 21981
rect 14553 22015 14611 22021
rect 14553 21981 14565 22015
rect 14599 22012 14611 22015
rect 14642 22012 14648 22024
rect 14599 21984 14648 22012
rect 14599 21981 14611 21984
rect 14553 21975 14611 21981
rect 14642 21972 14648 21984
rect 14700 21972 14706 22024
rect 14918 21972 14924 22024
rect 14976 22012 14982 22024
rect 15381 22015 15439 22021
rect 15381 22012 15393 22015
rect 14976 21984 15393 22012
rect 14976 21972 14982 21984
rect 15381 21981 15393 21984
rect 15427 21981 15439 22015
rect 15381 21975 15439 21981
rect 16574 21972 16580 22024
rect 16632 21972 16638 22024
rect 16684 21984 16896 22012
rect 6454 21904 6460 21956
rect 6512 21904 6518 21956
rect 6638 21904 6644 21956
rect 6696 21904 6702 21956
rect 16393 21947 16451 21953
rect 16393 21913 16405 21947
rect 16439 21944 16451 21947
rect 16684 21944 16712 21984
rect 16439 21916 16712 21944
rect 16439 21913 16451 21916
rect 16393 21907 16451 21913
rect 16758 21904 16764 21956
rect 16816 21904 16822 21956
rect 16868 21944 16896 21984
rect 17218 21972 17224 22024
rect 17276 21972 17282 22024
rect 17770 21972 17776 22024
rect 17828 22012 17834 22024
rect 18049 22015 18107 22021
rect 18049 22012 18061 22015
rect 17828 21984 18061 22012
rect 17828 21972 17834 21984
rect 18049 21981 18061 21984
rect 18095 21981 18107 22015
rect 18049 21975 18107 21981
rect 23658 21972 23664 22024
rect 23716 21972 23722 22024
rect 17313 21947 17371 21953
rect 17313 21944 17325 21947
rect 16868 21916 17325 21944
rect 17313 21913 17325 21916
rect 17359 21913 17371 21947
rect 17313 21907 17371 21913
rect 6822 21836 6828 21888
rect 6880 21836 6886 21888
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 12069 21879 12127 21885
rect 12069 21876 12081 21879
rect 12032 21848 12081 21876
rect 12032 21836 12038 21848
rect 12069 21845 12081 21848
rect 12115 21845 12127 21879
rect 12069 21839 12127 21845
rect 12529 21879 12587 21885
rect 12529 21845 12541 21879
rect 12575 21876 12587 21879
rect 12943 21879 13001 21885
rect 12943 21876 12955 21879
rect 12575 21848 12955 21876
rect 12575 21845 12587 21848
rect 12529 21839 12587 21845
rect 12943 21845 12955 21848
rect 12989 21845 13001 21879
rect 12943 21839 13001 21845
rect 14182 21836 14188 21888
rect 14240 21836 14246 21888
rect 14645 21879 14703 21885
rect 14645 21845 14657 21879
rect 14691 21876 14703 21879
rect 14734 21876 14740 21888
rect 14691 21848 14740 21876
rect 14691 21845 14703 21848
rect 14645 21839 14703 21845
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 16666 21836 16672 21888
rect 16724 21876 16730 21888
rect 16853 21879 16911 21885
rect 16853 21876 16865 21879
rect 16724 21848 16865 21876
rect 16724 21836 16730 21848
rect 16853 21845 16865 21848
rect 16899 21845 16911 21879
rect 16853 21839 16911 21845
rect 23477 21879 23535 21885
rect 23477 21845 23489 21879
rect 23523 21876 23535 21879
rect 23566 21876 23572 21888
rect 23523 21848 23572 21876
rect 23523 21845 23535 21848
rect 23477 21839 23535 21845
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 1104 21786 24012 21808
rect 1104 21734 4473 21786
rect 4525 21734 4537 21786
rect 4589 21734 4601 21786
rect 4653 21734 4665 21786
rect 4717 21734 4729 21786
rect 4781 21734 10200 21786
rect 10252 21734 10264 21786
rect 10316 21734 10328 21786
rect 10380 21734 10392 21786
rect 10444 21734 10456 21786
rect 10508 21734 15927 21786
rect 15979 21734 15991 21786
rect 16043 21734 16055 21786
rect 16107 21734 16119 21786
rect 16171 21734 16183 21786
rect 16235 21734 21654 21786
rect 21706 21734 21718 21786
rect 21770 21734 21782 21786
rect 21834 21734 21846 21786
rect 21898 21734 21910 21786
rect 21962 21734 24012 21786
rect 1104 21712 24012 21734
rect 1581 21675 1639 21681
rect 1581 21641 1593 21675
rect 1627 21672 1639 21675
rect 1627 21644 2774 21672
rect 1627 21641 1639 21644
rect 1581 21635 1639 21641
rect 842 21496 848 21548
rect 900 21536 906 21548
rect 1397 21539 1455 21545
rect 1397 21536 1409 21539
rect 900 21508 1409 21536
rect 900 21496 906 21508
rect 1397 21505 1409 21508
rect 1443 21505 1455 21539
rect 2746 21536 2774 21644
rect 3973 21607 4031 21613
rect 3973 21604 3985 21607
rect 3344 21576 3985 21604
rect 3344 21545 3372 21576
rect 3973 21573 3985 21576
rect 4019 21573 4031 21607
rect 3973 21567 4031 21573
rect 9861 21607 9919 21613
rect 9861 21573 9873 21607
rect 9907 21604 9919 21607
rect 9950 21604 9956 21616
rect 9907 21576 9956 21604
rect 9907 21573 9919 21576
rect 9861 21567 9919 21573
rect 9950 21564 9956 21576
rect 10008 21564 10014 21616
rect 15102 21604 15108 21616
rect 14752 21576 15108 21604
rect 3344 21539 3422 21545
rect 3344 21536 3376 21539
rect 2746 21508 3376 21536
rect 1397 21499 1455 21505
rect 3364 21505 3376 21508
rect 3410 21505 3422 21539
rect 3364 21499 3422 21505
rect 3467 21539 3525 21545
rect 3467 21505 3479 21539
rect 3513 21536 3525 21539
rect 3881 21539 3939 21545
rect 3881 21536 3893 21539
rect 3513 21508 3893 21536
rect 3513 21505 3525 21508
rect 3467 21499 3525 21505
rect 3881 21505 3893 21508
rect 3927 21505 3939 21539
rect 3881 21499 3939 21505
rect 4522 21496 4528 21548
rect 4580 21545 4586 21548
rect 4580 21539 4608 21545
rect 4596 21505 4608 21539
rect 4580 21499 4608 21505
rect 4580 21496 4586 21499
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 9125 21539 9183 21545
rect 9125 21536 9137 21539
rect 8996 21508 9137 21536
rect 8996 21496 9002 21508
rect 9125 21505 9137 21508
rect 9171 21536 9183 21539
rect 9214 21536 9220 21548
rect 9171 21508 9220 21536
rect 9171 21505 9183 21508
rect 9125 21499 9183 21505
rect 9214 21496 9220 21508
rect 9272 21496 9278 21548
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21536 9367 21539
rect 9677 21539 9735 21545
rect 9677 21536 9689 21539
rect 9355 21508 9689 21536
rect 9355 21505 9367 21508
rect 9309 21499 9367 21505
rect 9677 21505 9689 21508
rect 9723 21505 9735 21539
rect 11974 21536 11980 21548
rect 9677 21499 9735 21505
rect 11900 21508 11980 21536
rect 3789 21471 3847 21477
rect 3789 21437 3801 21471
rect 3835 21468 3847 21471
rect 5534 21468 5540 21480
rect 3835 21440 5540 21468
rect 3835 21437 3847 21440
rect 3789 21431 3847 21437
rect 5534 21428 5540 21440
rect 5592 21428 5598 21480
rect 6086 21428 6092 21480
rect 6144 21468 6150 21480
rect 6638 21468 6644 21480
rect 6144 21440 6644 21468
rect 6144 21428 6150 21440
rect 6638 21428 6644 21440
rect 6696 21468 6702 21480
rect 6733 21471 6791 21477
rect 6733 21468 6745 21471
rect 6696 21440 6745 21468
rect 6696 21428 6702 21440
rect 6733 21437 6745 21440
rect 6779 21468 6791 21471
rect 7193 21471 7251 21477
rect 7193 21468 7205 21471
rect 6779 21440 7205 21468
rect 6779 21437 6791 21440
rect 6733 21431 6791 21437
rect 7193 21437 7205 21440
rect 7239 21437 7251 21471
rect 7193 21431 7251 21437
rect 11238 21428 11244 21480
rect 11296 21468 11302 21480
rect 11900 21477 11928 21508
rect 11974 21496 11980 21508
rect 12032 21536 12038 21548
rect 14752 21545 14780 21576
rect 15102 21564 15108 21576
rect 15160 21564 15166 21616
rect 12345 21539 12403 21545
rect 12345 21536 12357 21539
rect 12032 21508 12357 21536
rect 12032 21496 12038 21508
rect 12345 21505 12357 21508
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 12529 21539 12587 21545
rect 12529 21505 12541 21539
rect 12575 21505 12587 21539
rect 12529 21499 12587 21505
rect 14737 21539 14795 21545
rect 14737 21505 14749 21539
rect 14783 21505 14795 21539
rect 14737 21499 14795 21505
rect 14921 21539 14979 21545
rect 14921 21505 14933 21539
rect 14967 21536 14979 21539
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 14967 21508 15301 21536
rect 14967 21505 14979 21508
rect 14921 21499 14979 21505
rect 15289 21505 15301 21508
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 15473 21499 15531 21505
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 11296 21440 11897 21468
rect 11296 21428 11302 21440
rect 11885 21437 11897 21440
rect 11931 21437 11943 21471
rect 12544 21468 12572 21499
rect 11885 21431 11943 21437
rect 12406 21440 12572 21468
rect 5994 21360 6000 21412
rect 6052 21400 6058 21412
rect 6454 21400 6460 21412
rect 6052 21372 6460 21400
rect 6052 21360 6058 21372
rect 6454 21360 6460 21372
rect 6512 21400 6518 21412
rect 6549 21403 6607 21409
rect 6549 21400 6561 21403
rect 6512 21372 6561 21400
rect 6512 21360 6518 21372
rect 6549 21369 6561 21372
rect 6595 21400 6607 21403
rect 7009 21403 7067 21409
rect 7009 21400 7021 21403
rect 6595 21372 7021 21400
rect 6595 21369 6607 21372
rect 6549 21363 6607 21369
rect 7009 21369 7021 21372
rect 7055 21369 7067 21403
rect 7009 21363 7067 21369
rect 8938 21360 8944 21412
rect 8996 21360 9002 21412
rect 12066 21360 12072 21412
rect 12124 21400 12130 21412
rect 12406 21400 12434 21440
rect 15102 21428 15108 21480
rect 15160 21468 15166 21480
rect 15488 21468 15516 21499
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17460 21508 17509 21536
rect 17460 21496 17466 21508
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21536 17739 21539
rect 17865 21539 17923 21545
rect 17865 21536 17877 21539
rect 17727 21508 17877 21536
rect 17727 21505 17739 21508
rect 17681 21499 17739 21505
rect 17865 21505 17877 21508
rect 17911 21505 17923 21539
rect 17865 21499 17923 21505
rect 18046 21496 18052 21548
rect 18104 21496 18110 21548
rect 18233 21539 18291 21545
rect 18233 21505 18245 21539
rect 18279 21536 18291 21539
rect 19613 21539 19671 21545
rect 19613 21536 19625 21539
rect 18279 21508 19625 21536
rect 18279 21505 18291 21508
rect 18233 21499 18291 21505
rect 19613 21505 19625 21508
rect 19659 21536 19671 21539
rect 23477 21539 23535 21545
rect 19659 21508 20116 21536
rect 19659 21505 19671 21508
rect 19613 21499 19671 21505
rect 15160 21440 15516 21468
rect 15160 21428 15166 21440
rect 16758 21428 16764 21480
rect 16816 21468 16822 21480
rect 17313 21471 17371 21477
rect 17313 21468 17325 21471
rect 16816 21440 17325 21468
rect 16816 21428 16822 21440
rect 17313 21437 17325 21440
rect 17359 21468 17371 21471
rect 17770 21468 17776 21480
rect 17359 21440 17776 21468
rect 17359 21437 17371 21440
rect 17313 21431 17371 21437
rect 17770 21428 17776 21440
rect 17828 21428 17834 21480
rect 19705 21471 19763 21477
rect 19705 21437 19717 21471
rect 19751 21468 19763 21471
rect 19886 21468 19892 21480
rect 19751 21440 19892 21468
rect 19751 21437 19763 21440
rect 19705 21431 19763 21437
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 20088 21477 20116 21508
rect 23477 21505 23489 21539
rect 23523 21536 23535 21539
rect 23750 21536 23756 21548
rect 23523 21508 23756 21536
rect 23523 21505 23535 21508
rect 23477 21499 23535 21505
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 20073 21471 20131 21477
rect 20073 21437 20085 21471
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21437 20315 21471
rect 20257 21431 20315 21437
rect 12124 21372 12434 21400
rect 14553 21403 14611 21409
rect 12124 21360 12130 21372
rect 14553 21369 14565 21403
rect 14599 21400 14611 21403
rect 14918 21400 14924 21412
rect 14599 21372 14924 21400
rect 14599 21369 14611 21372
rect 14553 21363 14611 21369
rect 14918 21360 14924 21372
rect 14976 21360 14982 21412
rect 19904 21400 19932 21428
rect 20272 21400 20300 21431
rect 20714 21428 20720 21480
rect 20772 21428 20778 21480
rect 20898 21428 20904 21480
rect 20956 21428 20962 21480
rect 19904 21372 20300 21400
rect 20441 21403 20499 21409
rect 20441 21369 20453 21403
rect 20487 21400 20499 21403
rect 20806 21400 20812 21412
rect 20487 21372 20812 21400
rect 20487 21369 20499 21372
rect 20441 21363 20499 21369
rect 20806 21360 20812 21372
rect 20864 21360 20870 21412
rect 4338 21292 4344 21344
rect 4396 21292 4402 21344
rect 4430 21292 4436 21344
rect 4488 21341 4494 21344
rect 4488 21335 4537 21341
rect 4488 21301 4491 21335
rect 4525 21301 4537 21335
rect 4488 21295 4537 21301
rect 6917 21335 6975 21341
rect 6917 21301 6929 21335
rect 6963 21332 6975 21335
rect 7282 21332 7288 21344
rect 6963 21304 7288 21332
rect 6963 21301 6975 21304
rect 6917 21295 6975 21301
rect 4488 21292 4494 21295
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7374 21292 7380 21344
rect 7432 21292 7438 21344
rect 9493 21335 9551 21341
rect 9493 21301 9505 21335
rect 9539 21332 9551 21335
rect 10318 21332 10324 21344
rect 9539 21304 10324 21332
rect 9539 21301 9551 21304
rect 9493 21295 9551 21301
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 11701 21335 11759 21341
rect 11701 21301 11713 21335
rect 11747 21332 11759 21335
rect 11790 21332 11796 21344
rect 11747 21304 11796 21332
rect 11747 21301 11759 21304
rect 11701 21295 11759 21301
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 11882 21292 11888 21344
rect 11940 21332 11946 21344
rect 12161 21335 12219 21341
rect 12161 21332 12173 21335
rect 11940 21304 12173 21332
rect 11940 21292 11946 21304
rect 12161 21301 12173 21304
rect 12207 21301 12219 21335
rect 12161 21295 12219 21301
rect 15657 21335 15715 21341
rect 15657 21301 15669 21335
rect 15703 21332 15715 21335
rect 16942 21332 16948 21344
rect 15703 21304 16948 21332
rect 15703 21301 15715 21304
rect 15657 21295 15715 21301
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 19794 21292 19800 21344
rect 19852 21332 19858 21344
rect 19981 21335 20039 21341
rect 19981 21332 19993 21335
rect 19852 21304 19993 21332
rect 19852 21292 19858 21304
rect 19981 21301 19993 21304
rect 20027 21301 20039 21335
rect 19981 21295 20039 21301
rect 20530 21292 20536 21344
rect 20588 21292 20594 21344
rect 23658 21292 23664 21344
rect 23716 21292 23722 21344
rect 1104 21242 24012 21264
rect 1104 21190 3813 21242
rect 3865 21190 3877 21242
rect 3929 21190 3941 21242
rect 3993 21190 4005 21242
rect 4057 21190 4069 21242
rect 4121 21190 9540 21242
rect 9592 21190 9604 21242
rect 9656 21190 9668 21242
rect 9720 21190 9732 21242
rect 9784 21190 9796 21242
rect 9848 21190 15267 21242
rect 15319 21190 15331 21242
rect 15383 21190 15395 21242
rect 15447 21190 15459 21242
rect 15511 21190 15523 21242
rect 15575 21190 20994 21242
rect 21046 21190 21058 21242
rect 21110 21190 21122 21242
rect 21174 21190 21186 21242
rect 21238 21190 21250 21242
rect 21302 21190 24012 21242
rect 1104 21168 24012 21190
rect 10318 21088 10324 21140
rect 10376 21128 10382 21140
rect 10376 21100 12756 21128
rect 10376 21088 10382 21100
rect 12728 21069 12756 21100
rect 15102 21088 15108 21140
rect 15160 21088 15166 21140
rect 17773 21131 17831 21137
rect 17773 21097 17785 21131
rect 17819 21128 17831 21131
rect 18046 21128 18052 21140
rect 17819 21100 18052 21128
rect 17819 21097 17831 21100
rect 17773 21091 17831 21097
rect 18046 21088 18052 21100
rect 18104 21088 18110 21140
rect 10781 21063 10839 21069
rect 10781 21060 10793 21063
rect 10428 21032 10793 21060
rect 4430 20952 4436 21004
rect 4488 20952 4494 21004
rect 4617 20995 4675 21001
rect 4617 20961 4629 20995
rect 4663 20992 4675 20995
rect 5902 20992 5908 21004
rect 4663 20964 5908 20992
rect 4663 20961 4675 20964
rect 4617 20955 4675 20961
rect 5902 20952 5908 20964
rect 5960 20952 5966 21004
rect 6086 20952 6092 21004
rect 6144 20952 6150 21004
rect 6362 20952 6368 21004
rect 6420 20952 6426 21004
rect 6822 20952 6828 21004
rect 6880 20992 6886 21004
rect 6917 20995 6975 21001
rect 6917 20992 6929 20995
rect 6880 20964 6929 20992
rect 6880 20952 6886 20964
rect 6917 20961 6929 20964
rect 6963 20961 6975 20995
rect 6917 20955 6975 20961
rect 7006 20952 7012 21004
rect 7064 20952 7070 21004
rect 9214 20952 9220 21004
rect 9272 20952 9278 21004
rect 9490 20952 9496 21004
rect 9548 20952 9554 21004
rect 10428 21001 10456 21032
rect 10781 21029 10793 21032
rect 10827 21060 10839 21063
rect 12713 21063 12771 21069
rect 10827 21032 12434 21060
rect 10827 21029 10839 21032
rect 10781 21023 10839 21029
rect 10413 20995 10471 21001
rect 10413 20961 10425 20995
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 10686 20952 10692 21004
rect 10744 20952 10750 21004
rect 11238 20952 11244 21004
rect 11296 20952 11302 21004
rect 11882 20952 11888 21004
rect 11940 20952 11946 21004
rect 12069 20995 12127 21001
rect 12069 20961 12081 20995
rect 12115 20992 12127 20995
rect 12158 20992 12164 21004
rect 12115 20964 12164 20992
rect 12115 20961 12127 20964
rect 12069 20955 12127 20961
rect 12158 20952 12164 20964
rect 12216 20952 12222 21004
rect 12253 20995 12311 21001
rect 12253 20961 12265 20995
rect 12299 20961 12311 20995
rect 12406 20992 12434 21032
rect 12713 21029 12725 21063
rect 12759 21029 12771 21063
rect 12713 21023 12771 21029
rect 17052 21032 17632 21060
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12406 20964 12909 20992
rect 12253 20955 12311 20961
rect 12897 20961 12909 20964
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 5994 20884 6000 20936
rect 6052 20884 6058 20936
rect 7282 20884 7288 20936
rect 7340 20884 7346 20936
rect 7653 20927 7711 20933
rect 7653 20893 7665 20927
rect 7699 20924 7711 20927
rect 8938 20924 8944 20936
rect 7699 20896 8944 20924
rect 7699 20893 7711 20896
rect 7653 20887 7711 20893
rect 8938 20884 8944 20896
rect 8996 20924 9002 20936
rect 9125 20927 9183 20933
rect 9125 20924 9137 20927
rect 8996 20896 9137 20924
rect 8996 20884 9002 20896
rect 9125 20893 9137 20896
rect 9171 20893 9183 20927
rect 9125 20887 9183 20893
rect 10318 20884 10324 20936
rect 10376 20884 10382 20936
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20924 11207 20927
rect 11195 20896 11744 20924
rect 11195 20893 11207 20896
rect 11149 20887 11207 20893
rect 4341 20859 4399 20865
rect 4341 20856 4353 20859
rect 2746 20828 4353 20856
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20788 1639 20791
rect 2746 20788 2774 20828
rect 4341 20825 4353 20828
rect 4387 20856 4399 20859
rect 4522 20856 4528 20868
rect 4387 20828 4528 20856
rect 4387 20825 4399 20828
rect 4341 20819 4399 20825
rect 4522 20816 4528 20828
rect 4580 20816 4586 20868
rect 6825 20859 6883 20865
rect 6825 20825 6837 20859
rect 6871 20856 6883 20859
rect 7374 20856 7380 20868
rect 6871 20828 7380 20856
rect 6871 20825 6883 20828
rect 6825 20819 6883 20825
rect 7374 20816 7380 20828
rect 7432 20816 7438 20868
rect 7466 20816 7472 20868
rect 7524 20816 7530 20868
rect 11238 20816 11244 20868
rect 11296 20856 11302 20868
rect 11716 20856 11744 20896
rect 11790 20884 11796 20936
rect 11848 20884 11854 20936
rect 12066 20856 12072 20868
rect 11296 20828 11560 20856
rect 11716 20828 12072 20856
rect 11296 20816 11302 20828
rect 1627 20760 2774 20788
rect 1627 20757 1639 20760
rect 1581 20751 1639 20757
rect 3694 20748 3700 20800
rect 3752 20788 3758 20800
rect 3973 20791 4031 20797
rect 3973 20788 3985 20791
rect 3752 20760 3985 20788
rect 3752 20748 3758 20760
rect 3973 20757 3985 20760
rect 4019 20757 4031 20791
rect 3973 20751 4031 20757
rect 6457 20791 6515 20797
rect 6457 20757 6469 20791
rect 6503 20788 6515 20791
rect 6730 20788 6736 20800
rect 6503 20760 6736 20788
rect 6503 20757 6515 20760
rect 6457 20751 6515 20757
rect 6730 20748 6736 20760
rect 6788 20748 6794 20800
rect 11422 20748 11428 20800
rect 11480 20748 11486 20800
rect 11532 20788 11560 20828
rect 12066 20816 12072 20828
rect 12124 20856 12130 20868
rect 12268 20856 12296 20955
rect 14734 20952 14740 21004
rect 14792 20952 14798 21004
rect 17052 21001 17080 21032
rect 17604 21004 17632 21032
rect 18138 21020 18144 21072
rect 18196 21060 18202 21072
rect 18196 21032 20024 21060
rect 18196 21020 18202 21032
rect 17037 20995 17095 21001
rect 17037 20961 17049 20995
rect 17083 20961 17095 20995
rect 17037 20955 17095 20961
rect 17310 20952 17316 21004
rect 17368 20952 17374 21004
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20961 17463 20995
rect 17405 20955 17463 20961
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20893 12495 20927
rect 12437 20887 12495 20893
rect 12452 20856 12480 20887
rect 14642 20884 14648 20936
rect 14700 20924 14706 20936
rect 14921 20927 14979 20933
rect 14921 20924 14933 20927
rect 14700 20896 14933 20924
rect 14700 20884 14706 20896
rect 14921 20893 14933 20896
rect 14967 20924 14979 20927
rect 15010 20924 15016 20936
rect 14967 20896 15016 20924
rect 14967 20893 14979 20896
rect 14921 20887 14979 20893
rect 15010 20884 15016 20896
rect 15068 20884 15074 20936
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17420 20924 17448 20955
rect 17586 20952 17592 21004
rect 17644 20952 17650 21004
rect 19996 21001 20024 21032
rect 20898 21020 20904 21072
rect 20956 21060 20962 21072
rect 21085 21063 21143 21069
rect 21085 21060 21097 21063
rect 20956 21032 21097 21060
rect 20956 21020 20962 21032
rect 21085 21029 21097 21032
rect 21131 21029 21143 21063
rect 21085 21023 21143 21029
rect 19061 20995 19119 21001
rect 19061 20961 19073 20995
rect 19107 20992 19119 20995
rect 19889 20995 19947 21001
rect 19889 20992 19901 20995
rect 19107 20964 19901 20992
rect 19107 20961 19119 20964
rect 19061 20955 19119 20961
rect 19889 20961 19901 20964
rect 19935 20961 19947 20995
rect 19889 20955 19947 20961
rect 19981 20995 20039 21001
rect 19981 20961 19993 20995
rect 20027 20992 20039 20995
rect 20809 20995 20867 21001
rect 20809 20992 20821 20995
rect 20027 20964 20821 20992
rect 20027 20961 20039 20964
rect 19981 20955 20039 20961
rect 20809 20961 20821 20964
rect 20855 20961 20867 20995
rect 20809 20955 20867 20961
rect 22738 20952 22744 21004
rect 22796 20952 22802 21004
rect 17000 20896 17448 20924
rect 17000 20884 17006 20896
rect 19794 20884 19800 20936
rect 19852 20884 19858 20936
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 21266 20924 21272 20936
rect 20772 20896 21272 20924
rect 20772 20884 20778 20896
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 23106 20933 23112 20936
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20924 22523 20927
rect 23074 20927 23112 20933
rect 23074 20924 23086 20927
rect 22511 20896 23086 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 23074 20893 23086 20896
rect 23074 20887 23112 20893
rect 23106 20884 23112 20887
rect 23164 20884 23170 20936
rect 23382 20884 23388 20936
rect 23440 20924 23446 20936
rect 23661 20927 23719 20933
rect 23661 20924 23673 20927
rect 23440 20896 23673 20924
rect 23440 20884 23446 20896
rect 23661 20893 23673 20896
rect 23707 20893 23719 20927
rect 23661 20887 23719 20893
rect 12124 20828 12296 20856
rect 12406 20828 12480 20856
rect 20625 20859 20683 20865
rect 12124 20816 12130 20828
rect 12406 20788 12434 20828
rect 20625 20825 20637 20859
rect 20671 20856 20683 20859
rect 21453 20859 21511 20865
rect 21453 20856 21465 20859
rect 20671 20828 21465 20856
rect 20671 20825 20683 20828
rect 20625 20819 20683 20825
rect 21453 20825 21465 20828
rect 21499 20825 21511 20859
rect 21453 20819 21511 20825
rect 11532 20760 12434 20788
rect 12618 20748 12624 20800
rect 12676 20748 12682 20800
rect 13078 20748 13084 20800
rect 13136 20748 13142 20800
rect 19426 20748 19432 20800
rect 19484 20748 19490 20800
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 20257 20791 20315 20797
rect 20257 20788 20269 20791
rect 19576 20760 20269 20788
rect 19576 20748 19582 20760
rect 20257 20757 20269 20760
rect 20303 20757 20315 20791
rect 20257 20751 20315 20757
rect 20714 20748 20720 20800
rect 20772 20748 20778 20800
rect 21266 20748 21272 20800
rect 21324 20788 21330 20800
rect 22097 20791 22155 20797
rect 22097 20788 22109 20791
rect 21324 20760 22109 20788
rect 21324 20748 21330 20760
rect 22097 20757 22109 20760
rect 22143 20757 22155 20791
rect 22097 20751 22155 20757
rect 22557 20791 22615 20797
rect 22557 20757 22569 20791
rect 22603 20788 22615 20791
rect 22971 20791 23029 20797
rect 22971 20788 22983 20791
rect 22603 20760 22983 20788
rect 22603 20757 22615 20760
rect 22557 20751 22615 20757
rect 22971 20757 22983 20760
rect 23017 20757 23029 20791
rect 22971 20751 23029 20757
rect 23474 20748 23480 20800
rect 23532 20748 23538 20800
rect 1104 20698 24012 20720
rect 1104 20646 4473 20698
rect 4525 20646 4537 20698
rect 4589 20646 4601 20698
rect 4653 20646 4665 20698
rect 4717 20646 4729 20698
rect 4781 20646 10200 20698
rect 10252 20646 10264 20698
rect 10316 20646 10328 20698
rect 10380 20646 10392 20698
rect 10444 20646 10456 20698
rect 10508 20646 15927 20698
rect 15979 20646 15991 20698
rect 16043 20646 16055 20698
rect 16107 20646 16119 20698
rect 16171 20646 16183 20698
rect 16235 20646 21654 20698
rect 21706 20646 21718 20698
rect 21770 20646 21782 20698
rect 21834 20646 21846 20698
rect 21898 20646 21910 20698
rect 21962 20646 24012 20698
rect 1104 20624 24012 20646
rect 6917 20587 6975 20593
rect 6917 20553 6929 20587
rect 6963 20584 6975 20587
rect 7466 20584 7472 20596
rect 6963 20556 7472 20584
rect 6963 20553 6975 20556
rect 6917 20547 6975 20553
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 9125 20587 9183 20593
rect 9125 20553 9137 20587
rect 9171 20584 9183 20587
rect 9490 20584 9496 20596
rect 9171 20556 9496 20584
rect 9171 20553 9183 20556
rect 9125 20547 9183 20553
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 14182 20544 14188 20596
rect 14240 20544 14246 20596
rect 17221 20587 17279 20593
rect 17221 20553 17233 20587
rect 17267 20584 17279 20587
rect 17310 20584 17316 20596
rect 17267 20556 17316 20584
rect 17267 20553 17279 20556
rect 17221 20547 17279 20553
rect 17310 20544 17316 20556
rect 17368 20544 17374 20596
rect 19426 20544 19432 20596
rect 19484 20544 19490 20596
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20772 20556 21005 20584
rect 20772 20544 20778 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 20993 20547 21051 20553
rect 12253 20519 12311 20525
rect 3712 20488 4108 20516
rect 3712 20460 3740 20488
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20448 3663 20451
rect 3694 20448 3700 20460
rect 3651 20420 3700 20448
rect 3651 20417 3663 20420
rect 3605 20411 3663 20417
rect 3694 20408 3700 20420
rect 3752 20408 3758 20460
rect 4080 20457 4108 20488
rect 12253 20485 12265 20519
rect 12299 20516 12311 20519
rect 12618 20516 12624 20528
rect 12299 20488 12624 20516
rect 12299 20485 12311 20488
rect 12253 20479 12311 20485
rect 12618 20476 12624 20488
rect 12676 20476 12682 20528
rect 19337 20519 19395 20525
rect 19337 20485 19349 20519
rect 19383 20516 19395 20519
rect 19518 20516 19524 20528
rect 19383 20488 19524 20516
rect 19383 20485 19395 20488
rect 19337 20479 19395 20485
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 20530 20476 20536 20528
rect 20588 20476 20594 20528
rect 20898 20516 20904 20528
rect 20640 20488 20904 20516
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20448 3847 20451
rect 4065 20451 4123 20457
rect 3835 20420 3924 20448
rect 3835 20417 3847 20420
rect 3789 20411 3847 20417
rect 3896 20321 3924 20420
rect 4065 20417 4077 20451
rect 4111 20448 4123 20451
rect 4525 20451 4583 20457
rect 4525 20448 4537 20451
rect 4111 20420 4537 20448
rect 4111 20417 4123 20420
rect 4065 20411 4123 20417
rect 4525 20417 4537 20420
rect 4571 20417 4583 20451
rect 4525 20411 4583 20417
rect 6362 20408 6368 20460
rect 6420 20448 6426 20460
rect 6733 20451 6791 20457
rect 6733 20448 6745 20451
rect 6420 20420 6745 20448
rect 6420 20408 6426 20420
rect 6733 20417 6745 20420
rect 6779 20417 6791 20451
rect 6733 20411 6791 20417
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9585 20451 9643 20457
rect 9585 20448 9597 20451
rect 9263 20420 9597 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 9585 20417 9597 20420
rect 9631 20417 9643 20451
rect 9585 20411 9643 20417
rect 12069 20451 12127 20457
rect 12069 20417 12081 20451
rect 12115 20417 12127 20451
rect 13078 20448 13084 20460
rect 12069 20411 12127 20417
rect 12406 20420 13084 20448
rect 4338 20340 4344 20392
rect 4396 20340 4402 20392
rect 9398 20340 9404 20392
rect 9456 20340 9462 20392
rect 12084 20380 12112 20411
rect 12406 20380 12434 20420
rect 13078 20408 13084 20420
rect 13136 20408 13142 20460
rect 14826 20448 14832 20460
rect 14016 20420 14832 20448
rect 14016 20389 14044 20420
rect 14826 20408 14832 20420
rect 14884 20408 14890 20460
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14976 20420 15025 20448
rect 14976 20408 14982 20420
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15013 20411 15071 20417
rect 15105 20451 15163 20457
rect 15105 20417 15117 20451
rect 15151 20448 15163 20451
rect 15473 20451 15531 20457
rect 15473 20448 15485 20451
rect 15151 20420 15485 20448
rect 15151 20417 15163 20420
rect 15105 20411 15163 20417
rect 15473 20417 15485 20420
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20448 17371 20451
rect 17681 20451 17739 20457
rect 17681 20448 17693 20451
rect 17359 20420 17693 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 17681 20417 17693 20420
rect 17727 20417 17739 20451
rect 17681 20411 17739 20417
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20448 20315 20451
rect 20640 20448 20668 20488
rect 20898 20476 20904 20488
rect 20956 20516 20962 20528
rect 21361 20519 21419 20525
rect 21361 20516 21373 20519
rect 20956 20488 21373 20516
rect 20956 20476 20962 20488
rect 21361 20485 21373 20488
rect 21407 20485 21419 20519
rect 21361 20479 21419 20485
rect 20303 20420 20668 20448
rect 20717 20451 20775 20457
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 20717 20417 20729 20451
rect 20763 20448 20775 20451
rect 20806 20448 20812 20460
rect 20763 20420 20812 20448
rect 20763 20417 20775 20420
rect 20717 20411 20775 20417
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 21177 20451 21235 20457
rect 21177 20417 21189 20451
rect 21223 20448 21235 20451
rect 21266 20448 21272 20460
rect 21223 20420 21272 20448
rect 21223 20417 21235 20420
rect 21177 20411 21235 20417
rect 12084 20352 12434 20380
rect 14001 20383 14059 20389
rect 14001 20349 14013 20383
rect 14047 20349 14059 20383
rect 14001 20343 14059 20349
rect 14093 20383 14151 20389
rect 14093 20349 14105 20383
rect 14139 20380 14151 20383
rect 15289 20383 15347 20389
rect 14139 20352 14688 20380
rect 14139 20349 14151 20352
rect 14093 20343 14151 20349
rect 3881 20315 3939 20321
rect 3881 20281 3893 20315
rect 3927 20312 3939 20315
rect 4356 20312 4384 20340
rect 3927 20284 4384 20312
rect 3927 20281 3939 20284
rect 3881 20275 3939 20281
rect 6546 20272 6552 20324
rect 6604 20272 6610 20324
rect 14660 20321 14688 20352
rect 15289 20349 15301 20383
rect 15335 20380 15347 20383
rect 17494 20380 17500 20392
rect 15335 20352 17500 20380
rect 15335 20349 15347 20352
rect 15289 20343 15347 20349
rect 17494 20340 17500 20352
rect 17552 20380 17558 20392
rect 17862 20380 17868 20392
rect 17552 20352 17868 20380
rect 17552 20340 17558 20352
rect 17862 20340 17868 20352
rect 17920 20340 17926 20392
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20380 19671 20383
rect 19794 20380 19800 20392
rect 19659 20352 19800 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 19794 20340 19800 20352
rect 19852 20340 19858 20392
rect 19886 20340 19892 20392
rect 19944 20340 19950 20392
rect 20349 20383 20407 20389
rect 20349 20349 20361 20383
rect 20395 20380 20407 20383
rect 21192 20380 21220 20411
rect 21266 20408 21272 20420
rect 21324 20408 21330 20460
rect 20395 20352 21220 20380
rect 20395 20349 20407 20352
rect 20349 20343 20407 20349
rect 14645 20315 14703 20321
rect 14645 20281 14657 20315
rect 14691 20281 14703 20315
rect 14645 20275 14703 20281
rect 3418 20204 3424 20256
rect 3476 20204 3482 20256
rect 4246 20204 4252 20256
rect 4304 20204 4310 20256
rect 4430 20204 4436 20256
rect 4488 20244 4494 20256
rect 4709 20247 4767 20253
rect 4709 20244 4721 20247
rect 4488 20216 4721 20244
rect 4488 20204 4494 20216
rect 4709 20213 4721 20216
rect 4755 20213 4767 20247
rect 4709 20207 4767 20213
rect 8757 20247 8815 20253
rect 8757 20213 8769 20247
rect 8803 20244 8815 20247
rect 8938 20244 8944 20256
rect 8803 20216 8944 20244
rect 8803 20213 8815 20216
rect 8757 20207 8815 20213
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 10594 20204 10600 20256
rect 10652 20204 10658 20256
rect 11885 20247 11943 20253
rect 11885 20213 11897 20247
rect 11931 20244 11943 20247
rect 12710 20244 12716 20256
rect 11931 20216 12716 20244
rect 11931 20213 11943 20216
rect 11885 20207 11943 20213
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 14090 20204 14096 20256
rect 14148 20244 14154 20256
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 14148 20216 14565 20244
rect 14148 20204 14154 20216
rect 14553 20213 14565 20216
rect 14599 20213 14611 20247
rect 14553 20207 14611 20213
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 16853 20247 16911 20253
rect 16853 20244 16865 20247
rect 16816 20216 16865 20244
rect 16816 20204 16822 20216
rect 16853 20213 16865 20216
rect 16899 20213 16911 20247
rect 16853 20207 16911 20213
rect 18966 20204 18972 20256
rect 19024 20204 19030 20256
rect 20898 20204 20904 20256
rect 20956 20204 20962 20256
rect 1104 20154 24012 20176
rect 1104 20102 3813 20154
rect 3865 20102 3877 20154
rect 3929 20102 3941 20154
rect 3993 20102 4005 20154
rect 4057 20102 4069 20154
rect 4121 20102 9540 20154
rect 9592 20102 9604 20154
rect 9656 20102 9668 20154
rect 9720 20102 9732 20154
rect 9784 20102 9796 20154
rect 9848 20102 15267 20154
rect 15319 20102 15331 20154
rect 15383 20102 15395 20154
rect 15447 20102 15459 20154
rect 15511 20102 15523 20154
rect 15575 20102 20994 20154
rect 21046 20102 21058 20154
rect 21110 20102 21122 20154
rect 21174 20102 21186 20154
rect 21238 20102 21250 20154
rect 21302 20102 24012 20154
rect 1104 20080 24012 20102
rect 14277 20043 14335 20049
rect 14277 20009 14289 20043
rect 14323 20040 14335 20043
rect 14458 20040 14464 20052
rect 14323 20012 14464 20040
rect 14323 20009 14335 20012
rect 14277 20003 14335 20009
rect 14458 20000 14464 20012
rect 14516 20000 14522 20052
rect 14918 20000 14924 20052
rect 14976 20000 14982 20052
rect 16025 20043 16083 20049
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 16390 20040 16396 20052
rect 16071 20012 16396 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 5350 19972 5356 19984
rect 4172 19944 5356 19972
rect 4172 19913 4200 19944
rect 5350 19932 5356 19944
rect 5408 19932 5414 19984
rect 9398 19932 9404 19984
rect 9456 19972 9462 19984
rect 9456 19944 10824 19972
rect 9456 19932 9462 19944
rect 4157 19907 4215 19913
rect 4157 19873 4169 19907
rect 4203 19873 4215 19907
rect 4157 19867 4215 19873
rect 4246 19864 4252 19916
rect 4304 19904 4310 19916
rect 4304 19876 4936 19904
rect 4304 19864 4310 19876
rect 842 19796 848 19848
rect 900 19836 906 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 900 19808 1409 19836
rect 900 19796 906 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 3418 19796 3424 19848
rect 3476 19836 3482 19848
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 3476 19808 4353 19836
rect 3476 19796 3482 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 4341 19799 4399 19805
rect 4430 19796 4436 19848
rect 4488 19796 4494 19848
rect 4908 19845 4936 19876
rect 6362 19864 6368 19916
rect 6420 19904 6426 19916
rect 6457 19907 6515 19913
rect 6457 19904 6469 19907
rect 6420 19876 6469 19904
rect 6420 19864 6426 19876
rect 6457 19873 6469 19876
rect 6503 19873 6515 19907
rect 6457 19867 6515 19873
rect 6914 19864 6920 19916
rect 6972 19864 6978 19916
rect 8754 19864 8760 19916
rect 8812 19904 8818 19916
rect 9861 19907 9919 19913
rect 9861 19904 9873 19907
rect 8812 19876 9873 19904
rect 8812 19864 8818 19876
rect 9861 19873 9873 19876
rect 9907 19873 9919 19907
rect 9861 19867 9919 19873
rect 10594 19864 10600 19916
rect 10652 19864 10658 19916
rect 10796 19913 10824 19944
rect 10781 19907 10839 19913
rect 10781 19873 10793 19907
rect 10827 19904 10839 19907
rect 12158 19904 12164 19916
rect 10827 19876 12164 19904
rect 10827 19873 10839 19876
rect 10781 19867 10839 19873
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 14642 19864 14648 19916
rect 14700 19864 14706 19916
rect 16758 19864 16764 19916
rect 16816 19864 16822 19916
rect 16942 19864 16948 19916
rect 17000 19864 17006 19916
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19805 4951 19839
rect 4893 19799 4951 19805
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19836 5319 19839
rect 6546 19836 6552 19848
rect 5307 19808 6552 19836
rect 5307 19805 5319 19808
rect 5261 19799 5319 19805
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 7009 19839 7067 19845
rect 7009 19805 7021 19839
rect 7055 19836 7067 19839
rect 7098 19836 7104 19848
rect 7055 19808 7104 19836
rect 7055 19805 7067 19808
rect 7009 19799 7067 19805
rect 7098 19796 7104 19808
rect 7156 19796 7162 19848
rect 9677 19839 9735 19845
rect 9677 19805 9689 19839
rect 9723 19836 9735 19839
rect 11422 19836 11428 19848
rect 9723 19808 11428 19836
rect 9723 19805 9735 19808
rect 9677 19799 9735 19805
rect 11422 19796 11428 19808
rect 11480 19796 11486 19848
rect 14090 19796 14096 19848
rect 14148 19796 14154 19848
rect 14553 19839 14611 19845
rect 14553 19805 14565 19839
rect 14599 19836 14611 19839
rect 14734 19836 14740 19848
rect 14599 19808 14740 19836
rect 14599 19805 14611 19808
rect 14553 19799 14611 19805
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 15838 19796 15844 19848
rect 15896 19796 15902 19848
rect 16666 19796 16672 19848
rect 16724 19796 16730 19848
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 23477 19839 23535 19845
rect 23477 19836 23489 19839
rect 18840 19808 23489 19836
rect 18840 19796 18846 19808
rect 23477 19805 23489 19808
rect 23523 19805 23535 19839
rect 23477 19799 23535 19805
rect 2593 19771 2651 19777
rect 2593 19737 2605 19771
rect 2639 19768 2651 19771
rect 4246 19768 4252 19780
rect 2639 19740 4252 19768
rect 2639 19737 2651 19740
rect 2593 19731 2651 19737
rect 4246 19728 4252 19740
rect 4304 19728 4310 19780
rect 5074 19728 5080 19780
rect 5132 19728 5138 19780
rect 10505 19771 10563 19777
rect 10505 19737 10517 19771
rect 10551 19768 10563 19771
rect 10686 19768 10692 19780
rect 10551 19740 10692 19768
rect 10551 19737 10563 19740
rect 10505 19731 10563 19737
rect 10686 19728 10692 19740
rect 10744 19728 10750 19780
rect 4798 19660 4804 19712
rect 4856 19660 4862 19712
rect 9309 19703 9367 19709
rect 9309 19669 9321 19703
rect 9355 19700 9367 19703
rect 9398 19700 9404 19712
rect 9355 19672 9404 19700
rect 9355 19669 9367 19672
rect 9309 19663 9367 19669
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 10137 19703 10195 19709
rect 10137 19700 10149 19703
rect 9815 19672 10149 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 10137 19669 10149 19672
rect 10183 19669 10195 19703
rect 10137 19663 10195 19669
rect 15838 19660 15844 19712
rect 15896 19700 15902 19712
rect 16301 19703 16359 19709
rect 16301 19700 16313 19703
rect 15896 19672 16313 19700
rect 15896 19660 15902 19672
rect 16301 19669 16313 19672
rect 16347 19669 16359 19703
rect 16301 19663 16359 19669
rect 23658 19660 23664 19712
rect 23716 19660 23722 19712
rect 1104 19610 24012 19632
rect 1104 19558 4473 19610
rect 4525 19558 4537 19610
rect 4589 19558 4601 19610
rect 4653 19558 4665 19610
rect 4717 19558 4729 19610
rect 4781 19558 10200 19610
rect 10252 19558 10264 19610
rect 10316 19558 10328 19610
rect 10380 19558 10392 19610
rect 10444 19558 10456 19610
rect 10508 19558 15927 19610
rect 15979 19558 15991 19610
rect 16043 19558 16055 19610
rect 16107 19558 16119 19610
rect 16171 19558 16183 19610
rect 16235 19558 21654 19610
rect 21706 19558 21718 19610
rect 21770 19558 21782 19610
rect 21834 19558 21846 19610
rect 21898 19558 21910 19610
rect 21962 19558 24012 19610
rect 1104 19536 24012 19558
rect 6914 19456 6920 19508
rect 6972 19496 6978 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 6972 19468 7021 19496
rect 6972 19456 6978 19468
rect 7009 19465 7021 19468
rect 7055 19465 7067 19499
rect 7009 19459 7067 19465
rect 7098 19456 7104 19508
rect 7156 19456 7162 19508
rect 8938 19456 8944 19508
rect 8996 19456 9002 19508
rect 9030 19456 9036 19508
rect 9088 19456 9094 19508
rect 18782 19456 18788 19508
rect 18840 19456 18846 19508
rect 23382 19456 23388 19508
rect 23440 19456 23446 19508
rect 23477 19499 23535 19505
rect 23477 19465 23489 19499
rect 23523 19496 23535 19499
rect 23658 19496 23664 19508
rect 23523 19468 23664 19496
rect 23523 19465 23535 19468
rect 23477 19459 23535 19465
rect 23658 19456 23664 19468
rect 23716 19456 23722 19508
rect 7190 19428 7196 19440
rect 2746 19400 7196 19428
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19360 1639 19363
rect 2746 19360 2774 19400
rect 7190 19388 7196 19400
rect 7248 19388 7254 19440
rect 1627 19332 2774 19360
rect 3789 19363 3847 19369
rect 1627 19329 1639 19332
rect 1581 19323 1639 19329
rect 3789 19329 3801 19363
rect 3835 19360 3847 19363
rect 4338 19360 4344 19372
rect 3835 19332 4344 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 14826 19360 14832 19372
rect 8772 19332 14832 19360
rect 8772 19304 8800 19332
rect 14826 19320 14832 19332
rect 14884 19360 14890 19372
rect 16942 19360 16948 19372
rect 14884 19332 16948 19360
rect 14884 19320 14890 19332
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 18230 19320 18236 19372
rect 18288 19360 18294 19372
rect 18601 19363 18659 19369
rect 18601 19360 18613 19363
rect 18288 19332 18613 19360
rect 18288 19320 18294 19332
rect 18601 19329 18613 19332
rect 18647 19360 18659 19363
rect 18966 19360 18972 19372
rect 18647 19332 18972 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 23198 19320 23204 19372
rect 23256 19320 23262 19372
rect 23290 19320 23296 19372
rect 23348 19360 23354 19372
rect 23661 19363 23719 19369
rect 23661 19360 23673 19363
rect 23348 19332 23673 19360
rect 23348 19320 23354 19332
rect 23661 19329 23673 19332
rect 23707 19329 23719 19363
rect 23661 19323 23719 19329
rect 3694 19252 3700 19304
rect 3752 19252 3758 19304
rect 7006 19252 7012 19304
rect 7064 19292 7070 19304
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 7064 19264 7297 19292
rect 7064 19252 7070 19264
rect 7285 19261 7297 19264
rect 7331 19292 7343 19295
rect 8202 19292 8208 19304
rect 7331 19264 8208 19292
rect 7331 19261 7343 19264
rect 7285 19255 7343 19261
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 8754 19252 8760 19304
rect 8812 19252 8818 19304
rect 1394 19116 1400 19168
rect 1452 19116 1458 19168
rect 4154 19116 4160 19168
rect 4212 19116 4218 19168
rect 6638 19116 6644 19168
rect 6696 19116 6702 19168
rect 8938 19116 8944 19168
rect 8996 19156 9002 19168
rect 9401 19159 9459 19165
rect 9401 19156 9413 19159
rect 8996 19128 9413 19156
rect 8996 19116 9002 19128
rect 9401 19125 9413 19128
rect 9447 19125 9459 19159
rect 9401 19119 9459 19125
rect 1104 19066 24012 19088
rect 1104 19014 3813 19066
rect 3865 19014 3877 19066
rect 3929 19014 3941 19066
rect 3993 19014 4005 19066
rect 4057 19014 4069 19066
rect 4121 19014 9540 19066
rect 9592 19014 9604 19066
rect 9656 19014 9668 19066
rect 9720 19014 9732 19066
rect 9784 19014 9796 19066
rect 9848 19014 15267 19066
rect 15319 19014 15331 19066
rect 15383 19014 15395 19066
rect 15447 19014 15459 19066
rect 15511 19014 15523 19066
rect 15575 19014 20994 19066
rect 21046 19014 21058 19066
rect 21110 19014 21122 19066
rect 21174 19014 21186 19066
rect 21238 19014 21250 19066
rect 21302 19014 24012 19066
rect 1104 18992 24012 19014
rect 4157 18955 4215 18961
rect 4157 18921 4169 18955
rect 4203 18952 4215 18955
rect 5074 18952 5080 18964
rect 4203 18924 5080 18952
rect 4203 18921 4215 18924
rect 4157 18915 4215 18921
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 7190 18912 7196 18964
rect 7248 18912 7254 18964
rect 9122 18912 9128 18964
rect 9180 18912 9186 18964
rect 9585 18955 9643 18961
rect 9585 18921 9597 18955
rect 9631 18952 9643 18955
rect 10042 18952 10048 18964
rect 9631 18924 10048 18952
rect 9631 18921 9643 18924
rect 9585 18915 9643 18921
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 14369 18955 14427 18961
rect 14369 18921 14381 18955
rect 14415 18952 14427 18955
rect 15838 18952 15844 18964
rect 14415 18924 15844 18952
rect 14415 18921 14427 18924
rect 14369 18915 14427 18921
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 18325 18955 18383 18961
rect 18325 18921 18337 18955
rect 18371 18952 18383 18955
rect 23198 18952 23204 18964
rect 18371 18924 23204 18952
rect 18371 18921 18383 18924
rect 18325 18915 18383 18921
rect 23198 18912 23204 18924
rect 23256 18912 23262 18964
rect 12636 18856 13216 18884
rect 12636 18828 12664 18856
rect 3789 18819 3847 18825
rect 3789 18785 3801 18819
rect 3835 18816 3847 18819
rect 4246 18816 4252 18828
rect 3835 18788 4252 18816
rect 3835 18785 3847 18788
rect 3789 18779 3847 18785
rect 4246 18776 4252 18788
rect 4304 18776 4310 18828
rect 4430 18776 4436 18828
rect 4488 18816 4494 18828
rect 4890 18816 4896 18828
rect 4488 18788 4896 18816
rect 4488 18776 4494 18788
rect 4890 18776 4896 18788
rect 4948 18816 4954 18828
rect 6457 18819 6515 18825
rect 6457 18816 6469 18819
rect 4948 18788 6469 18816
rect 4948 18776 4954 18788
rect 6457 18785 6469 18788
rect 6503 18785 6515 18819
rect 6457 18779 6515 18785
rect 6638 18776 6644 18828
rect 6696 18776 6702 18828
rect 12158 18776 12164 18828
rect 12216 18776 12222 18828
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 1627 18720 2774 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 2746 18680 2774 18720
rect 3970 18708 3976 18760
rect 4028 18708 4034 18760
rect 4617 18751 4675 18757
rect 4617 18717 4629 18751
rect 4663 18748 4675 18751
rect 4798 18748 4804 18760
rect 4663 18720 4804 18748
rect 4663 18717 4675 18720
rect 4617 18711 4675 18717
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 5074 18708 5080 18760
rect 5132 18708 5138 18760
rect 6730 18708 6736 18760
rect 6788 18708 6794 18760
rect 7377 18751 7435 18757
rect 7377 18748 7389 18751
rect 7116 18720 7389 18748
rect 7006 18680 7012 18692
rect 2746 18652 7012 18680
rect 7006 18640 7012 18652
rect 7064 18640 7070 18692
rect 7116 18624 7144 18720
rect 7377 18717 7389 18720
rect 7423 18717 7435 18751
rect 7377 18711 7435 18717
rect 8938 18708 8944 18760
rect 8996 18708 9002 18760
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 11885 18751 11943 18757
rect 11885 18717 11897 18751
rect 11931 18748 11943 18751
rect 12360 18748 12388 18779
rect 12618 18776 12624 18828
rect 12676 18776 12682 18828
rect 13188 18825 13216 18856
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 14645 18887 14703 18893
rect 14148 18856 14504 18884
rect 14148 18844 14154 18856
rect 14476 18825 14504 18856
rect 14645 18853 14657 18887
rect 14691 18884 14703 18887
rect 14734 18884 14740 18896
rect 14691 18856 14740 18884
rect 14691 18853 14703 18856
rect 14645 18847 14703 18853
rect 14734 18844 14740 18856
rect 14792 18844 14798 18896
rect 12989 18819 13047 18825
rect 12989 18785 13001 18819
rect 13035 18785 13047 18819
rect 12989 18779 13047 18785
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18785 13231 18819
rect 13173 18779 13231 18785
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18785 14335 18819
rect 14277 18779 14335 18785
rect 14461 18819 14519 18825
rect 14461 18785 14473 18819
rect 14507 18785 14519 18819
rect 14461 18779 14519 18785
rect 11931 18720 12388 18748
rect 11931 18717 11943 18720
rect 11885 18711 11943 18717
rect 12710 18708 12716 18760
rect 12768 18748 12774 18760
rect 13004 18748 13032 18779
rect 12768 18720 13032 18748
rect 14292 18748 14320 18779
rect 19794 18776 19800 18828
rect 19852 18776 19858 18828
rect 21913 18819 21971 18825
rect 21913 18816 21925 18819
rect 19904 18788 21925 18816
rect 17681 18751 17739 18757
rect 14292 18720 17632 18748
rect 12768 18708 12774 18720
rect 14090 18640 14096 18692
rect 14148 18640 14154 18692
rect 14550 18640 14556 18692
rect 14608 18680 14614 18692
rect 14829 18683 14887 18689
rect 14829 18680 14841 18683
rect 14608 18652 14841 18680
rect 14608 18640 14614 18652
rect 14829 18649 14841 18652
rect 14875 18649 14887 18683
rect 14829 18643 14887 18649
rect 15013 18683 15071 18689
rect 15013 18649 15025 18683
rect 15059 18680 15071 18683
rect 15286 18680 15292 18692
rect 15059 18652 15292 18680
rect 15059 18649 15071 18652
rect 15013 18643 15071 18649
rect 15286 18640 15292 18652
rect 15344 18640 15350 18692
rect 17604 18680 17632 18720
rect 17681 18717 17693 18751
rect 17727 18748 17739 18751
rect 18046 18748 18052 18760
rect 17727 18720 18052 18748
rect 17727 18717 17739 18720
rect 17681 18711 17739 18717
rect 18046 18708 18052 18720
rect 18104 18708 18110 18760
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 18156 18680 18184 18711
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19904 18748 19932 18788
rect 21913 18785 21925 18788
rect 21959 18785 21971 18819
rect 21913 18779 21971 18785
rect 23014 18776 23020 18828
rect 23072 18816 23078 18828
rect 23198 18816 23204 18828
rect 23072 18788 23204 18816
rect 23072 18776 23078 18788
rect 23198 18776 23204 18788
rect 23256 18776 23262 18828
rect 19300 18720 19932 18748
rect 19300 18708 19306 18720
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 20073 18751 20131 18757
rect 20073 18748 20085 18751
rect 20036 18720 20085 18748
rect 20036 18708 20042 18720
rect 20073 18717 20085 18720
rect 20119 18717 20131 18751
rect 20073 18711 20131 18717
rect 22925 18751 22983 18757
rect 22925 18717 22937 18751
rect 22971 18748 22983 18751
rect 23474 18748 23480 18760
rect 23532 18757 23538 18760
rect 23532 18751 23560 18757
rect 22971 18720 23480 18748
rect 22971 18717 22983 18720
rect 22925 18711 22983 18717
rect 23474 18708 23480 18720
rect 23548 18717 23560 18751
rect 23532 18711 23560 18717
rect 23532 18708 23538 18711
rect 19613 18683 19671 18689
rect 17604 18652 19288 18680
rect 842 18572 848 18624
rect 900 18612 906 18624
rect 1397 18615 1455 18621
rect 1397 18612 1409 18615
rect 900 18584 1409 18612
rect 900 18572 906 18584
rect 1397 18581 1409 18584
rect 1443 18581 1455 18615
rect 1397 18575 1455 18581
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 4525 18615 4583 18621
rect 4525 18612 4537 18615
rect 4304 18584 4537 18612
rect 4304 18572 4310 18584
rect 4525 18581 4537 18584
rect 4571 18581 4583 18615
rect 4525 18575 4583 18581
rect 4982 18572 4988 18624
rect 5040 18572 5046 18624
rect 7098 18572 7104 18624
rect 7156 18572 7162 18624
rect 11514 18572 11520 18624
rect 11572 18572 11578 18624
rect 11974 18572 11980 18624
rect 12032 18572 12038 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 13357 18615 13415 18621
rect 13357 18612 13369 18615
rect 13320 18584 13369 18612
rect 13320 18572 13326 18584
rect 13357 18581 13369 18584
rect 13403 18581 13415 18615
rect 13357 18575 13415 18581
rect 13998 18572 14004 18624
rect 14056 18612 14062 18624
rect 19260 18621 19288 18652
rect 19613 18649 19625 18683
rect 19659 18680 19671 18683
rect 21729 18683 21787 18689
rect 19659 18652 21404 18680
rect 19659 18649 19671 18652
rect 19613 18643 19671 18649
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 14056 18584 14197 18612
rect 14056 18572 14062 18584
rect 14185 18581 14197 18584
rect 14231 18581 14243 18615
rect 14185 18575 14243 18581
rect 19245 18615 19303 18621
rect 19245 18581 19257 18615
rect 19291 18581 19303 18615
rect 19245 18575 19303 18581
rect 19518 18572 19524 18624
rect 19576 18612 19582 18624
rect 21376 18621 21404 18652
rect 21729 18649 21741 18683
rect 21775 18680 21787 18683
rect 22094 18680 22100 18692
rect 21775 18652 22100 18680
rect 21775 18649 21787 18652
rect 21729 18643 21787 18649
rect 22094 18640 22100 18652
rect 22152 18640 22158 18692
rect 19705 18615 19763 18621
rect 19705 18612 19717 18615
rect 19576 18584 19717 18612
rect 19576 18572 19582 18584
rect 19705 18581 19717 18584
rect 19751 18581 19763 18615
rect 19705 18575 19763 18581
rect 21361 18615 21419 18621
rect 21361 18581 21373 18615
rect 21407 18581 21419 18615
rect 21361 18575 21419 18581
rect 21821 18615 21879 18621
rect 21821 18581 21833 18615
rect 21867 18612 21879 18615
rect 22370 18612 22376 18624
rect 21867 18584 22376 18612
rect 21867 18581 21879 18584
rect 21821 18575 21879 18581
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 22554 18572 22560 18624
rect 22612 18572 22618 18624
rect 23017 18615 23075 18621
rect 23017 18581 23029 18615
rect 23063 18612 23075 18615
rect 23431 18615 23489 18621
rect 23431 18612 23443 18615
rect 23063 18584 23443 18612
rect 23063 18581 23075 18584
rect 23017 18575 23075 18581
rect 23431 18581 23443 18584
rect 23477 18581 23489 18615
rect 23431 18575 23489 18581
rect 1104 18522 24012 18544
rect 1104 18470 4473 18522
rect 4525 18470 4537 18522
rect 4589 18470 4601 18522
rect 4653 18470 4665 18522
rect 4717 18470 4729 18522
rect 4781 18470 10200 18522
rect 10252 18470 10264 18522
rect 10316 18470 10328 18522
rect 10380 18470 10392 18522
rect 10444 18470 10456 18522
rect 10508 18470 15927 18522
rect 15979 18470 15991 18522
rect 16043 18470 16055 18522
rect 16107 18470 16119 18522
rect 16171 18470 16183 18522
rect 16235 18470 21654 18522
rect 21706 18470 21718 18522
rect 21770 18470 21782 18522
rect 21834 18470 21846 18522
rect 21898 18470 21910 18522
rect 21962 18470 24012 18522
rect 1104 18448 24012 18470
rect 4246 18368 4252 18420
rect 4304 18368 4310 18420
rect 4709 18411 4767 18417
rect 4709 18377 4721 18411
rect 4755 18408 4767 18411
rect 5074 18408 5080 18420
rect 4755 18380 5080 18408
rect 4755 18377 4767 18380
rect 4709 18371 4767 18377
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 8662 18368 8668 18420
rect 8720 18408 8726 18420
rect 8849 18411 8907 18417
rect 8849 18408 8861 18411
rect 8720 18380 8861 18408
rect 8720 18368 8726 18380
rect 8849 18377 8861 18380
rect 8895 18377 8907 18411
rect 8849 18371 8907 18377
rect 14550 18368 14556 18420
rect 14608 18368 14614 18420
rect 15286 18368 15292 18420
rect 15344 18368 15350 18420
rect 17221 18411 17279 18417
rect 17221 18377 17233 18411
rect 17267 18408 17279 18411
rect 17773 18411 17831 18417
rect 17773 18408 17785 18411
rect 17267 18380 17785 18408
rect 17267 18377 17279 18380
rect 17221 18371 17279 18377
rect 17773 18377 17785 18380
rect 17819 18377 17831 18411
rect 17773 18371 17831 18377
rect 18046 18368 18052 18420
rect 18104 18408 18110 18420
rect 18233 18411 18291 18417
rect 18233 18408 18245 18411
rect 18104 18380 18245 18408
rect 18104 18368 18110 18380
rect 18233 18377 18245 18380
rect 18279 18377 18291 18411
rect 18233 18371 18291 18377
rect 19518 18368 19524 18420
rect 19576 18368 19582 18420
rect 19978 18368 19984 18420
rect 20036 18368 20042 18420
rect 4338 18340 4344 18352
rect 3804 18312 4344 18340
rect 3804 18281 3832 18312
rect 4338 18300 4344 18312
rect 4396 18300 4402 18352
rect 9398 18300 9404 18352
rect 9456 18340 9462 18352
rect 9493 18343 9551 18349
rect 9493 18340 9505 18343
rect 9456 18312 9505 18340
rect 9456 18300 9462 18312
rect 9493 18309 9505 18312
rect 9539 18309 9551 18343
rect 9493 18303 9551 18309
rect 13262 18300 13268 18352
rect 13320 18300 13326 18352
rect 18141 18343 18199 18349
rect 18141 18340 18153 18343
rect 15212 18312 18153 18340
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 3789 18275 3847 18281
rect 1627 18244 2774 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 2746 18136 2774 18244
rect 3789 18241 3801 18275
rect 3835 18241 3847 18275
rect 4617 18275 4675 18281
rect 4617 18272 4629 18275
rect 3789 18235 3847 18241
rect 4172 18244 4629 18272
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18204 3939 18207
rect 3970 18204 3976 18216
rect 3927 18176 3976 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 4172 18213 4200 18244
rect 4617 18241 4629 18244
rect 4663 18241 4675 18275
rect 4617 18235 4675 18241
rect 4982 18232 4988 18284
rect 5040 18272 5046 18284
rect 9033 18275 9091 18281
rect 9033 18272 9045 18275
rect 5040 18244 9045 18272
rect 5040 18232 5046 18244
rect 9033 18241 9045 18244
rect 9079 18272 9091 18275
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 9079 18244 9229 18272
rect 9079 18241 9091 18244
rect 9033 18235 9091 18241
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18272 11943 18275
rect 11974 18272 11980 18284
rect 11931 18244 11980 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 11974 18232 11980 18244
rect 12032 18232 12038 18284
rect 13078 18232 13084 18284
rect 13136 18232 13142 18284
rect 14829 18275 14887 18281
rect 14829 18241 14841 18275
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18173 4215 18207
rect 4157 18167 4215 18173
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 5350 18204 5356 18216
rect 4939 18176 5356 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 9125 18207 9183 18213
rect 9125 18173 9137 18207
rect 9171 18204 9183 18207
rect 9398 18204 9404 18216
rect 9171 18176 9404 18204
rect 9171 18173 9183 18176
rect 9125 18167 9183 18173
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 14369 18207 14427 18213
rect 14369 18173 14381 18207
rect 14415 18204 14427 18207
rect 14734 18204 14740 18216
rect 14415 18176 14740 18204
rect 14415 18173 14427 18176
rect 14369 18167 14427 18173
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 6086 18136 6092 18148
rect 2746 18108 6092 18136
rect 6086 18096 6092 18108
rect 6144 18096 6150 18148
rect 8938 18096 8944 18148
rect 8996 18136 9002 18148
rect 9309 18139 9367 18145
rect 9309 18136 9321 18139
rect 8996 18108 9321 18136
rect 8996 18096 9002 18108
rect 9309 18105 9321 18108
rect 9355 18105 9367 18139
rect 9309 18099 9367 18105
rect 9493 18139 9551 18145
rect 9493 18105 9505 18139
rect 9539 18136 9551 18139
rect 13449 18139 13507 18145
rect 9539 18108 12434 18136
rect 9539 18105 9551 18108
rect 9493 18099 9551 18105
rect 1394 18028 1400 18080
rect 1452 18028 1458 18080
rect 12406 18068 12434 18108
rect 13449 18105 13461 18139
rect 13495 18136 13507 18139
rect 14185 18139 14243 18145
rect 14185 18136 14197 18139
rect 13495 18108 14197 18136
rect 13495 18105 13507 18108
rect 13449 18099 13507 18105
rect 14185 18105 14197 18108
rect 14231 18136 14243 18139
rect 14844 18136 14872 18235
rect 15212 18213 15240 18312
rect 18141 18309 18153 18312
rect 18187 18309 18199 18343
rect 18141 18303 18199 18309
rect 22925 18343 22983 18349
rect 22925 18309 22937 18343
rect 22971 18340 22983 18343
rect 22971 18312 23612 18340
rect 22971 18309 22983 18312
rect 22925 18303 22983 18309
rect 23584 18284 23612 18312
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15672 18244 15761 18272
rect 15197 18207 15255 18213
rect 15197 18173 15209 18207
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 14231 18108 14872 18136
rect 14231 18105 14243 18108
rect 14185 18099 14243 18105
rect 13170 18068 13176 18080
rect 12406 18040 13176 18068
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 15488 18068 15516 18167
rect 15672 18148 15700 18244
rect 15749 18241 15761 18244
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15896 18244 15945 18272
rect 15896 18232 15902 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 17310 18232 17316 18284
rect 17368 18232 17374 18284
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18272 19947 18275
rect 20717 18275 20775 18281
rect 19935 18244 20392 18272
rect 19935 18241 19947 18244
rect 19889 18235 19947 18241
rect 16942 18164 16948 18216
rect 17000 18204 17006 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 17000 18176 17141 18204
rect 17000 18164 17006 18176
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17129 18167 17187 18173
rect 15654 18096 15660 18148
rect 15712 18096 15718 18148
rect 17144 18136 17172 18167
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 18196 18176 18337 18204
rect 18196 18164 18202 18176
rect 18325 18173 18337 18176
rect 18371 18204 18383 18207
rect 19242 18204 19248 18216
rect 18371 18176 19248 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 19242 18164 19248 18176
rect 19300 18204 19306 18216
rect 20364 18213 20392 18244
rect 20717 18241 20729 18275
rect 20763 18272 20775 18275
rect 20898 18272 20904 18284
rect 20763 18244 20904 18272
rect 20763 18241 20775 18244
rect 20717 18235 20775 18241
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18272 22247 18275
rect 22554 18272 22560 18284
rect 22235 18244 22560 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 23566 18281 23572 18284
rect 23017 18275 23075 18281
rect 23017 18241 23029 18275
rect 23063 18272 23075 18275
rect 23431 18275 23489 18281
rect 23431 18272 23443 18275
rect 23063 18244 23443 18272
rect 23063 18241 23075 18244
rect 23017 18235 23075 18241
rect 23431 18241 23443 18244
rect 23477 18241 23489 18275
rect 23431 18235 23489 18241
rect 23534 18275 23572 18281
rect 23534 18241 23546 18275
rect 23534 18235 23572 18241
rect 23566 18232 23572 18235
rect 23624 18232 23630 18284
rect 20073 18207 20131 18213
rect 20073 18204 20085 18207
rect 19300 18176 20085 18204
rect 19300 18164 19306 18176
rect 20073 18173 20085 18176
rect 20119 18173 20131 18207
rect 20073 18167 20131 18173
rect 20349 18207 20407 18213
rect 20349 18173 20361 18207
rect 20395 18173 20407 18207
rect 20349 18167 20407 18173
rect 20809 18207 20867 18213
rect 20809 18173 20821 18207
rect 20855 18173 20867 18207
rect 20916 18204 20944 18232
rect 20993 18207 21051 18213
rect 20993 18204 21005 18207
rect 20916 18176 21005 18204
rect 20809 18167 20867 18173
rect 20993 18173 21005 18176
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 21177 18207 21235 18213
rect 21177 18173 21189 18207
rect 21223 18204 21235 18207
rect 21821 18207 21879 18213
rect 21821 18204 21833 18207
rect 21223 18176 21833 18204
rect 21223 18173 21235 18176
rect 21177 18167 21235 18173
rect 21821 18173 21833 18176
rect 21867 18173 21879 18207
rect 21821 18167 21879 18173
rect 22097 18207 22155 18213
rect 22097 18173 22109 18207
rect 22143 18173 22155 18207
rect 22097 18167 22155 18173
rect 19794 18136 19800 18148
rect 17144 18108 19800 18136
rect 19794 18096 19800 18108
rect 19852 18096 19858 18148
rect 20824 18136 20852 18167
rect 21192 18136 21220 18167
rect 20824 18108 21220 18136
rect 22112 18136 22140 18167
rect 22738 18164 22744 18216
rect 22796 18204 22802 18216
rect 23106 18204 23112 18216
rect 22796 18176 23112 18204
rect 22796 18164 22802 18176
rect 23106 18164 23112 18176
rect 23164 18164 23170 18216
rect 22278 18136 22284 18148
rect 22112 18108 22284 18136
rect 22278 18096 22284 18108
rect 22336 18136 22342 18148
rect 22557 18139 22615 18145
rect 22557 18136 22569 18139
rect 22336 18108 22569 18136
rect 22336 18096 22342 18108
rect 22557 18105 22569 18108
rect 22603 18105 22615 18139
rect 22557 18099 22615 18105
rect 15838 18068 15844 18080
rect 15488 18040 15844 18068
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 16117 18071 16175 18077
rect 16117 18037 16129 18071
rect 16163 18068 16175 18071
rect 16574 18068 16580 18080
rect 16163 18040 16580 18068
rect 16163 18037 16175 18040
rect 16117 18031 16175 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 17681 18071 17739 18077
rect 17681 18037 17693 18071
rect 17727 18068 17739 18071
rect 17862 18068 17868 18080
rect 17727 18040 17868 18068
rect 17727 18037 17739 18040
rect 17681 18031 17739 18037
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 21358 18028 21364 18080
rect 21416 18028 21422 18080
rect 1104 17978 24012 18000
rect 1104 17926 3813 17978
rect 3865 17926 3877 17978
rect 3929 17926 3941 17978
rect 3993 17926 4005 17978
rect 4057 17926 4069 17978
rect 4121 17926 9540 17978
rect 9592 17926 9604 17978
rect 9656 17926 9668 17978
rect 9720 17926 9732 17978
rect 9784 17926 9796 17978
rect 9848 17926 15267 17978
rect 15319 17926 15331 17978
rect 15383 17926 15395 17978
rect 15447 17926 15459 17978
rect 15511 17926 15523 17978
rect 15575 17926 20994 17978
rect 21046 17926 21058 17978
rect 21110 17926 21122 17978
rect 21174 17926 21186 17978
rect 21238 17926 21250 17978
rect 21302 17926 24012 17978
rect 1104 17904 24012 17926
rect 6086 17824 6092 17876
rect 6144 17824 6150 17876
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 7098 17864 7104 17876
rect 6595 17836 7104 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 9858 17824 9864 17876
rect 9916 17824 9922 17876
rect 12618 17824 12624 17876
rect 12676 17824 12682 17876
rect 13078 17824 13084 17876
rect 13136 17824 13142 17876
rect 14734 17824 14740 17876
rect 14792 17824 14798 17876
rect 16945 17867 17003 17873
rect 16945 17833 16957 17867
rect 16991 17864 17003 17867
rect 17310 17864 17316 17876
rect 16991 17836 17316 17864
rect 16991 17833 17003 17836
rect 16945 17827 17003 17833
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 22094 17824 22100 17876
rect 22152 17824 22158 17876
rect 22370 17824 22376 17876
rect 22428 17864 22434 17876
rect 22925 17867 22983 17873
rect 22925 17864 22937 17867
rect 22428 17836 22937 17864
rect 22428 17824 22434 17836
rect 22925 17833 22937 17836
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 6822 17796 6828 17808
rect 6380 17768 6828 17796
rect 6380 17737 6408 17768
rect 6822 17756 6828 17768
rect 6880 17756 6886 17808
rect 8754 17796 8760 17808
rect 7392 17768 8760 17796
rect 7392 17737 7420 17768
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 9585 17799 9643 17805
rect 9585 17765 9597 17799
rect 9631 17796 9643 17799
rect 11054 17796 11060 17808
rect 9631 17768 11060 17796
rect 9631 17765 9643 17768
rect 9585 17759 9643 17765
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 12713 17799 12771 17805
rect 12713 17796 12725 17799
rect 12268 17768 12725 17796
rect 6365 17731 6423 17737
rect 6365 17697 6377 17731
rect 6411 17697 6423 17731
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 6365 17691 6423 17697
rect 6656 17700 7389 17728
rect 6270 17620 6276 17672
rect 6328 17660 6334 17672
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 6328 17632 6469 17660
rect 6328 17620 6334 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 4798 17552 4804 17604
rect 4856 17592 4862 17604
rect 6656 17592 6684 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 8202 17688 8208 17740
rect 8260 17688 8266 17740
rect 8772 17728 8800 17756
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 8772 17700 10977 17728
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8481 17663 8539 17669
rect 8481 17660 8493 17663
rect 8159 17632 8493 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 8481 17629 8493 17632
rect 8527 17629 8539 17663
rect 8481 17623 8539 17629
rect 9398 17620 9404 17672
rect 9456 17620 9462 17672
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17660 10931 17663
rect 11514 17660 11520 17672
rect 10919 17632 11520 17660
rect 10919 17629 10931 17632
rect 10873 17623 10931 17629
rect 4856 17564 6684 17592
rect 6733 17595 6791 17601
rect 4856 17552 4862 17564
rect 6733 17561 6745 17595
rect 6779 17592 6791 17595
rect 9692 17592 9720 17623
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 12268 17669 12296 17768
rect 12713 17765 12725 17768
rect 12759 17765 12771 17799
rect 18138 17796 18144 17808
rect 12713 17759 12771 17765
rect 15028 17768 15884 17796
rect 15028 17737 15056 17768
rect 12345 17731 12403 17737
rect 12345 17697 12357 17731
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 15013 17731 15071 17737
rect 15013 17697 15025 17731
rect 15059 17697 15071 17731
rect 15013 17691 15071 17697
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17629 12311 17663
rect 12360 17660 12388 17691
rect 15654 17688 15660 17740
rect 15712 17688 15718 17740
rect 12618 17660 12624 17672
rect 12360 17632 12624 17660
rect 12253 17623 12311 17629
rect 12268 17592 12296 17623
rect 12618 17620 12624 17632
rect 12676 17660 12682 17672
rect 12897 17663 12955 17669
rect 12897 17660 12909 17663
rect 12676 17632 12909 17660
rect 12676 17620 12682 17632
rect 12897 17629 12909 17632
rect 12943 17629 12955 17663
rect 12897 17623 12955 17629
rect 15105 17663 15163 17669
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15194 17660 15200 17672
rect 15151 17632 15200 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 15194 17620 15200 17632
rect 15252 17660 15258 17672
rect 15672 17660 15700 17688
rect 15856 17672 15884 17768
rect 16408 17768 18144 17796
rect 16408 17737 16436 17768
rect 18138 17756 18144 17768
rect 18196 17756 18202 17808
rect 21177 17799 21235 17805
rect 21177 17765 21189 17799
rect 21223 17796 21235 17799
rect 22186 17796 22192 17808
rect 21223 17768 22192 17796
rect 21223 17765 21235 17768
rect 21177 17759 21235 17765
rect 22186 17756 22192 17768
rect 22244 17756 22250 17808
rect 22465 17799 22523 17805
rect 22465 17765 22477 17799
rect 22511 17796 22523 17799
rect 22554 17796 22560 17808
rect 22511 17768 22560 17796
rect 22511 17765 22523 17768
rect 22465 17759 22523 17765
rect 22554 17756 22560 17768
rect 22612 17756 22618 17808
rect 23658 17756 23664 17808
rect 23716 17756 23722 17808
rect 16393 17731 16451 17737
rect 16393 17697 16405 17731
rect 16439 17697 16451 17731
rect 16393 17691 16451 17697
rect 16485 17731 16543 17737
rect 16485 17697 16497 17731
rect 16531 17728 16543 17731
rect 16574 17728 16580 17740
rect 16531 17700 16580 17728
rect 16531 17697 16543 17700
rect 16485 17691 16543 17697
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22572 17728 22600 17756
rect 22051 17700 22600 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 15252 17632 15700 17660
rect 15252 17620 15258 17632
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 17862 17620 17868 17672
rect 17920 17620 17926 17672
rect 21358 17620 21364 17672
rect 21416 17620 21422 17672
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17660 21879 17663
rect 22278 17660 22284 17672
rect 21867 17632 22284 17660
rect 21867 17629 21879 17632
rect 21821 17623 21879 17629
rect 22278 17620 22284 17632
rect 22336 17620 22342 17672
rect 22572 17669 22600 17700
rect 22557 17663 22615 17669
rect 22557 17629 22569 17663
rect 22603 17629 22615 17663
rect 23477 17663 23535 17669
rect 23477 17660 23489 17663
rect 22557 17623 22615 17629
rect 22848 17632 23489 17660
rect 12342 17592 12348 17604
rect 6779 17564 10456 17592
rect 12268 17564 12348 17592
rect 6779 17561 6791 17564
rect 6733 17555 6791 17561
rect 6638 17484 6644 17536
rect 6696 17484 6702 17536
rect 7190 17484 7196 17536
rect 7248 17484 7254 17536
rect 7285 17527 7343 17533
rect 7285 17493 7297 17527
rect 7331 17524 7343 17527
rect 7653 17527 7711 17533
rect 7653 17524 7665 17527
rect 7331 17496 7665 17524
rect 7331 17493 7343 17496
rect 7285 17487 7343 17493
rect 7653 17493 7665 17496
rect 7699 17493 7711 17527
rect 7653 17487 7711 17493
rect 8018 17484 8024 17536
rect 8076 17484 8082 17536
rect 10428 17533 10456 17564
rect 12342 17552 12348 17564
rect 12400 17552 12406 17604
rect 16025 17595 16083 17601
rect 16025 17561 16037 17595
rect 16071 17592 16083 17595
rect 16577 17595 16635 17601
rect 16577 17592 16589 17595
rect 16071 17564 16589 17592
rect 16071 17561 16083 17564
rect 16025 17555 16083 17561
rect 16577 17561 16589 17564
rect 16623 17561 16635 17595
rect 21545 17595 21603 17601
rect 16577 17555 16635 17561
rect 18064 17564 21312 17592
rect 10413 17527 10471 17533
rect 10413 17493 10425 17527
rect 10459 17493 10471 17527
rect 10413 17487 10471 17493
rect 10778 17484 10784 17536
rect 10836 17484 10842 17536
rect 18064 17533 18092 17564
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17493 18107 17527
rect 21284 17524 21312 17564
rect 21545 17561 21557 17595
rect 21591 17592 21603 17595
rect 21637 17595 21695 17601
rect 21637 17592 21649 17595
rect 21591 17564 21649 17592
rect 21591 17561 21603 17564
rect 21545 17555 21603 17561
rect 21637 17561 21649 17564
rect 21683 17561 21695 17595
rect 22296 17592 22324 17620
rect 22741 17595 22799 17601
rect 22741 17592 22753 17595
rect 22296 17564 22753 17592
rect 21637 17555 21695 17561
rect 22741 17561 22753 17564
rect 22787 17561 22799 17595
rect 22741 17555 22799 17561
rect 22848 17524 22876 17632
rect 23477 17629 23489 17632
rect 23523 17629 23535 17663
rect 23477 17623 23535 17629
rect 21284 17496 22876 17524
rect 18049 17487 18107 17493
rect 1104 17434 24012 17456
rect 1104 17382 4473 17434
rect 4525 17382 4537 17434
rect 4589 17382 4601 17434
rect 4653 17382 4665 17434
rect 4717 17382 4729 17434
rect 4781 17382 10200 17434
rect 10252 17382 10264 17434
rect 10316 17382 10328 17434
rect 10380 17382 10392 17434
rect 10444 17382 10456 17434
rect 10508 17382 15927 17434
rect 15979 17382 15991 17434
rect 16043 17382 16055 17434
rect 16107 17382 16119 17434
rect 16171 17382 16183 17434
rect 16235 17382 21654 17434
rect 21706 17382 21718 17434
rect 21770 17382 21782 17434
rect 21834 17382 21846 17434
rect 21898 17382 21910 17434
rect 21962 17382 24012 17434
rect 1104 17360 24012 17382
rect 5353 17323 5411 17329
rect 5353 17289 5365 17323
rect 5399 17320 5411 17323
rect 6270 17320 6276 17332
rect 5399 17292 6276 17320
rect 5399 17289 5411 17292
rect 5353 17283 5411 17289
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 7006 17280 7012 17332
rect 7064 17280 7070 17332
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 10836 17292 11621 17320
rect 10836 17280 10842 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 15105 17323 15163 17329
rect 15105 17289 15117 17323
rect 15151 17320 15163 17323
rect 15194 17320 15200 17332
rect 15151 17292 15200 17320
rect 15151 17289 15163 17292
rect 15105 17283 15163 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 23566 17320 23572 17332
rect 16224 17292 23572 17320
rect 6638 17212 6644 17264
rect 6696 17252 6702 17264
rect 13538 17252 13544 17264
rect 6696 17224 13544 17252
rect 6696 17212 6702 17224
rect 13538 17212 13544 17224
rect 13596 17212 13602 17264
rect 15473 17255 15531 17261
rect 15473 17221 15485 17255
rect 15519 17252 15531 17255
rect 16224 17252 16252 17292
rect 23566 17280 23572 17292
rect 23624 17280 23630 17332
rect 15519 17224 16252 17252
rect 15519 17221 15531 17224
rect 15473 17215 15531 17221
rect 842 17144 848 17196
rect 900 17184 906 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 900 17156 1409 17184
rect 900 17144 906 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 4982 17144 4988 17196
rect 5040 17144 5046 17196
rect 6822 17144 6828 17196
rect 6880 17184 6886 17196
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6880 17156 7205 17184
rect 6880 17144 6886 17156
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17184 12035 17187
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12023 17156 12449 17184
rect 12023 17153 12035 17156
rect 11977 17147 12035 17153
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 12618 17144 12624 17196
rect 12676 17144 12682 17196
rect 12710 17144 12716 17196
rect 12768 17184 12774 17196
rect 13046 17187 13104 17193
rect 13046 17184 13058 17187
rect 12768 17156 13058 17184
rect 12768 17144 12774 17156
rect 13046 17153 13058 17156
rect 13092 17184 13104 17187
rect 13630 17184 13636 17196
rect 13092 17156 13636 17184
rect 13092 17153 13104 17156
rect 13046 17147 13104 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17184 15623 17187
rect 15979 17187 16037 17193
rect 15979 17184 15991 17187
rect 15611 17156 15991 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 15979 17153 15991 17156
rect 16025 17153 16037 17187
rect 15979 17147 16037 17153
rect 16082 17187 16140 17193
rect 16082 17153 16094 17187
rect 16128 17184 16140 17187
rect 16224 17184 16252 17224
rect 17862 17212 17868 17264
rect 17920 17252 17926 17264
rect 17957 17255 18015 17261
rect 17957 17252 17969 17255
rect 17920 17224 17969 17252
rect 17920 17212 17926 17224
rect 17957 17221 17969 17224
rect 18003 17221 18015 17255
rect 17957 17215 18015 17221
rect 18049 17187 18107 17193
rect 16128 17156 16252 17184
rect 16358 17179 16416 17185
rect 16128 17153 16140 17156
rect 16082 17147 16140 17153
rect 16358 17145 16370 17179
rect 16404 17145 16416 17179
rect 18049 17153 18061 17187
rect 18095 17184 18107 17187
rect 18230 17184 18236 17196
rect 18095 17156 18236 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 16358 17139 16416 17145
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17184 18935 17187
rect 19518 17184 19524 17196
rect 18923 17156 19524 17184
rect 18923 17153 18935 17156
rect 18877 17147 18935 17153
rect 4798 17076 4804 17128
rect 4856 17076 4862 17128
rect 4890 17076 4896 17128
rect 4948 17076 4954 17128
rect 12066 17076 12072 17128
rect 12124 17076 12130 17128
rect 12158 17076 12164 17128
rect 12216 17076 12222 17128
rect 13722 17076 13728 17128
rect 13780 17116 13786 17128
rect 15749 17119 15807 17125
rect 15749 17116 15761 17119
rect 13780 17088 15761 17116
rect 13780 17076 13786 17088
rect 15749 17085 15761 17088
rect 15795 17116 15807 17119
rect 16206 17116 16212 17128
rect 15795 17088 16212 17116
rect 15795 17085 15807 17088
rect 15749 17079 15807 17085
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 11790 17048 11796 17060
rect 2746 17020 11796 17048
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16980 1639 16983
rect 2746 16980 2774 17020
rect 11790 17008 11796 17020
rect 11848 17008 11854 17060
rect 12176 17048 12204 17076
rect 12084 17020 12204 17048
rect 1627 16952 2774 16980
rect 1627 16949 1639 16952
rect 1581 16943 1639 16949
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 11054 16940 11060 16992
rect 11112 16980 11118 16992
rect 12084 16980 12112 17020
rect 12342 17008 12348 17060
rect 12400 17048 12406 17060
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 12400 17020 12817 17048
rect 12400 17008 12406 17020
rect 12805 17017 12817 17020
rect 12851 17017 12863 17051
rect 12805 17011 12863 17017
rect 16114 17008 16120 17060
rect 16172 17048 16178 17060
rect 16383 17048 16411 17139
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17116 18199 17119
rect 18892 17116 18920 17147
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 23477 17187 23535 17193
rect 23477 17184 23489 17187
rect 22066 17156 23489 17184
rect 18187 17088 18920 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 19061 17051 19119 17057
rect 16172 17020 18460 17048
rect 16172 17008 16178 17020
rect 11112 16952 12112 16980
rect 11112 16940 11118 16952
rect 12894 16940 12900 16992
rect 12952 16989 12958 16992
rect 12952 16983 13001 16989
rect 12952 16949 12955 16983
rect 12989 16949 13001 16983
rect 12952 16943 13001 16949
rect 12952 16940 12958 16943
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16255 16983 16313 16989
rect 16255 16980 16267 16983
rect 15988 16952 16267 16980
rect 15988 16940 15994 16952
rect 16255 16949 16267 16952
rect 16301 16949 16313 16983
rect 16255 16943 16313 16949
rect 18230 16940 18236 16992
rect 18288 16980 18294 16992
rect 18325 16983 18383 16989
rect 18325 16980 18337 16983
rect 18288 16952 18337 16980
rect 18288 16940 18294 16952
rect 18325 16949 18337 16952
rect 18371 16949 18383 16983
rect 18432 16980 18460 17020
rect 19061 17017 19073 17051
rect 19107 17048 19119 17051
rect 22066 17048 22094 17156
rect 23477 17153 23489 17156
rect 23523 17153 23535 17187
rect 23477 17147 23535 17153
rect 19107 17020 22094 17048
rect 19107 17017 19119 17020
rect 19061 17011 19119 17017
rect 23658 17008 23664 17060
rect 23716 17008 23722 17060
rect 23842 16980 23848 16992
rect 18432 16952 23848 16980
rect 18325 16943 18383 16949
rect 23842 16940 23848 16952
rect 23900 16940 23906 16992
rect 1104 16890 24012 16912
rect 1104 16838 3813 16890
rect 3865 16838 3877 16890
rect 3929 16838 3941 16890
rect 3993 16838 4005 16890
rect 4057 16838 4069 16890
rect 4121 16838 9540 16890
rect 9592 16838 9604 16890
rect 9656 16838 9668 16890
rect 9720 16838 9732 16890
rect 9784 16838 9796 16890
rect 9848 16838 15267 16890
rect 15319 16838 15331 16890
rect 15383 16838 15395 16890
rect 15447 16838 15459 16890
rect 15511 16838 15523 16890
rect 15575 16838 20994 16890
rect 21046 16838 21058 16890
rect 21110 16838 21122 16890
rect 21174 16838 21186 16890
rect 21238 16838 21250 16890
rect 21302 16838 24012 16890
rect 1104 16816 24012 16838
rect 4801 16779 4859 16785
rect 4801 16745 4813 16779
rect 4847 16776 4859 16779
rect 4890 16776 4896 16788
rect 4847 16748 4896 16776
rect 4847 16745 4859 16748
rect 4801 16739 4859 16745
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 7101 16779 7159 16785
rect 7101 16745 7113 16779
rect 7147 16776 7159 16779
rect 7190 16776 7196 16788
rect 7147 16748 7196 16776
rect 7147 16745 7159 16748
rect 7101 16739 7159 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 9398 16736 9404 16788
rect 9456 16736 9462 16788
rect 11977 16779 12035 16785
rect 11977 16745 11989 16779
rect 12023 16776 12035 16779
rect 12066 16776 12072 16788
rect 12023 16748 12072 16776
rect 12023 16745 12035 16748
rect 11977 16739 12035 16745
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 12618 16776 12624 16788
rect 12483 16748 12624 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 5442 16708 5448 16720
rect 5276 16680 5448 16708
rect 5276 16649 5304 16680
rect 5442 16668 5448 16680
rect 5500 16668 5506 16720
rect 8202 16708 8208 16720
rect 7760 16680 8208 16708
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 5261 16603 5319 16609
rect 5350 16600 5356 16652
rect 5408 16640 5414 16652
rect 7760 16649 7788 16680
rect 8202 16668 8208 16680
rect 8260 16708 8266 16720
rect 11054 16708 11060 16720
rect 8260 16680 11060 16708
rect 8260 16668 8266 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 7745 16643 7803 16649
rect 7745 16640 7757 16643
rect 5408 16612 7757 16640
rect 5408 16600 5414 16612
rect 7745 16609 7757 16612
rect 7791 16609 7803 16643
rect 7745 16603 7803 16609
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 9953 16643 10011 16649
rect 9953 16640 9965 16643
rect 8904 16612 9965 16640
rect 8904 16600 8910 16612
rect 9953 16609 9965 16612
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 842 16532 848 16584
rect 900 16572 906 16584
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 900 16544 1409 16572
rect 900 16532 906 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 2746 16544 9996 16572
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16436 1639 16439
rect 2746 16436 2774 16544
rect 9766 16464 9772 16516
rect 9824 16464 9830 16516
rect 1627 16408 2774 16436
rect 1627 16405 1639 16408
rect 1581 16399 1639 16405
rect 5166 16396 5172 16448
rect 5224 16396 5230 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7469 16439 7527 16445
rect 7469 16436 7481 16439
rect 6972 16408 7481 16436
rect 6972 16396 6978 16408
rect 7469 16405 7481 16408
rect 7515 16405 7527 16439
rect 7469 16399 7527 16405
rect 7558 16396 7564 16448
rect 7616 16396 7622 16448
rect 9858 16396 9864 16448
rect 9916 16396 9922 16448
rect 9968 16436 9996 16544
rect 10042 16532 10048 16584
rect 10100 16572 10106 16584
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 10100 16544 10241 16572
rect 10100 16532 10106 16544
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 12342 16532 12348 16584
rect 12400 16532 12406 16584
rect 12161 16507 12219 16513
rect 12161 16473 12173 16507
rect 12207 16473 12219 16507
rect 12452 16504 12480 16739
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 15473 16779 15531 16785
rect 15473 16745 15485 16779
rect 15519 16776 15531 16779
rect 15838 16776 15844 16788
rect 15519 16748 15844 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 18322 16736 18328 16788
rect 18380 16776 18386 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 18380 16748 18429 16776
rect 18380 16736 18386 16748
rect 18417 16745 18429 16748
rect 18463 16745 18475 16779
rect 18417 16739 18475 16745
rect 19518 16736 19524 16788
rect 19576 16736 19582 16788
rect 13096 16680 16068 16708
rect 13096 16652 13124 16680
rect 13078 16600 13084 16652
rect 13136 16600 13142 16652
rect 15930 16600 15936 16652
rect 15988 16600 15994 16652
rect 16040 16649 16068 16680
rect 16206 16668 16212 16720
rect 16264 16708 16270 16720
rect 22002 16708 22008 16720
rect 16264 16680 22008 16708
rect 16264 16668 16270 16680
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 16025 16643 16083 16649
rect 16025 16609 16037 16643
rect 16071 16609 16083 16643
rect 16025 16603 16083 16609
rect 17865 16643 17923 16649
rect 17865 16609 17877 16643
rect 17911 16640 17923 16643
rect 18322 16640 18328 16652
rect 17911 16612 18328 16640
rect 17911 16609 17923 16612
rect 17865 16603 17923 16609
rect 18322 16600 18328 16612
rect 18380 16640 18386 16652
rect 19794 16640 19800 16652
rect 18380 16612 19800 16640
rect 18380 16600 18386 16612
rect 19794 16600 19800 16612
rect 19852 16640 19858 16652
rect 20073 16643 20131 16649
rect 20073 16640 20085 16643
rect 19852 16612 20085 16640
rect 19852 16600 19858 16612
rect 20073 16609 20085 16612
rect 20119 16609 20131 16643
rect 20073 16603 20131 16609
rect 12802 16532 12808 16584
rect 12860 16572 12866 16584
rect 13382 16575 13440 16581
rect 13382 16572 13394 16575
rect 12860 16544 13394 16572
rect 12860 16532 12866 16544
rect 13382 16541 13394 16544
rect 13428 16541 13440 16575
rect 13382 16535 13440 16541
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16572 15899 16575
rect 16114 16572 16120 16584
rect 15887 16544 16120 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 16114 16532 16120 16544
rect 16172 16532 16178 16584
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 18509 16575 18567 16581
rect 18509 16572 18521 16575
rect 18472 16544 18521 16572
rect 18472 16532 18478 16544
rect 18509 16541 18521 16544
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 18782 16532 18788 16584
rect 18840 16532 18846 16584
rect 20714 16532 20720 16584
rect 20772 16532 20778 16584
rect 23658 16532 23664 16584
rect 23716 16532 23722 16584
rect 23750 16504 23756 16516
rect 12161 16467 12219 16473
rect 12406 16476 12480 16504
rect 18708 16476 23756 16504
rect 11882 16436 11888 16448
rect 9968 16408 11888 16436
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 12176 16436 12204 16467
rect 12406 16436 12434 16476
rect 12176 16408 12434 16436
rect 12897 16439 12955 16445
rect 12897 16405 12909 16439
rect 12943 16436 12955 16439
rect 13311 16439 13369 16445
rect 13311 16436 13323 16439
rect 12943 16408 13323 16436
rect 12943 16405 12955 16408
rect 12897 16399 12955 16405
rect 13311 16405 13323 16408
rect 13357 16405 13369 16439
rect 13311 16399 13369 16405
rect 17954 16396 17960 16448
rect 18012 16396 18018 16448
rect 18046 16396 18052 16448
rect 18104 16396 18110 16448
rect 18708 16445 18736 16476
rect 23750 16464 23756 16476
rect 23808 16464 23814 16516
rect 18693 16439 18751 16445
rect 18693 16405 18705 16439
rect 18739 16405 18751 16439
rect 18693 16399 18751 16405
rect 19886 16396 19892 16448
rect 19944 16396 19950 16448
rect 19978 16396 19984 16448
rect 20036 16396 20042 16448
rect 23474 16396 23480 16448
rect 23532 16396 23538 16448
rect 1104 16346 24012 16368
rect 1104 16294 4473 16346
rect 4525 16294 4537 16346
rect 4589 16294 4601 16346
rect 4653 16294 4665 16346
rect 4717 16294 4729 16346
rect 4781 16294 10200 16346
rect 10252 16294 10264 16346
rect 10316 16294 10328 16346
rect 10380 16294 10392 16346
rect 10444 16294 10456 16346
rect 10508 16294 15927 16346
rect 15979 16294 15991 16346
rect 16043 16294 16055 16346
rect 16107 16294 16119 16346
rect 16171 16294 16183 16346
rect 16235 16294 21654 16346
rect 21706 16294 21718 16346
rect 21770 16294 21782 16346
rect 21834 16294 21846 16346
rect 21898 16294 21910 16346
rect 21962 16294 24012 16346
rect 1104 16272 24012 16294
rect 4338 16192 4344 16244
rect 4396 16192 4402 16244
rect 7377 16235 7435 16241
rect 7377 16201 7389 16235
rect 7423 16232 7435 16235
rect 7558 16232 7564 16244
rect 7423 16204 7564 16232
rect 7423 16201 7435 16204
rect 7377 16195 7435 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 9677 16235 9735 16241
rect 9677 16201 9689 16235
rect 9723 16232 9735 16235
rect 9858 16232 9864 16244
rect 9723 16204 9864 16232
rect 9723 16201 9735 16204
rect 9677 16195 9735 16201
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 10137 16235 10195 16241
rect 10137 16232 10149 16235
rect 10100 16204 10149 16232
rect 10100 16192 10106 16204
rect 10137 16201 10149 16204
rect 10183 16201 10195 16235
rect 10137 16195 10195 16201
rect 12342 16192 12348 16244
rect 12400 16192 12406 16244
rect 12710 16192 12716 16244
rect 12768 16192 12774 16244
rect 12805 16235 12863 16241
rect 12805 16201 12817 16235
rect 12851 16232 12863 16235
rect 12894 16232 12900 16244
rect 12851 16204 12900 16232
rect 12851 16201 12863 16204
rect 12805 16195 12863 16201
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 14277 16235 14335 16241
rect 14277 16201 14289 16235
rect 14323 16232 14335 16235
rect 15746 16232 15752 16244
rect 14323 16204 15752 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18141 16235 18199 16241
rect 18141 16232 18153 16235
rect 18012 16204 18153 16232
rect 18012 16192 18018 16204
rect 18141 16201 18153 16204
rect 18187 16201 18199 16235
rect 18141 16195 18199 16201
rect 18601 16235 18659 16241
rect 18601 16201 18613 16235
rect 18647 16232 18659 16235
rect 18782 16232 18788 16244
rect 18647 16204 18788 16232
rect 18647 16201 18659 16204
rect 18601 16195 18659 16201
rect 18782 16192 18788 16204
rect 18840 16192 18846 16244
rect 19978 16192 19984 16244
rect 20036 16232 20042 16244
rect 20349 16235 20407 16241
rect 20349 16232 20361 16235
rect 20036 16204 20361 16232
rect 20036 16192 20042 16204
rect 20349 16201 20361 16204
rect 20395 16201 20407 16235
rect 20349 16195 20407 16201
rect 20714 16192 20720 16244
rect 20772 16232 20778 16244
rect 20809 16235 20867 16241
rect 20809 16232 20821 16235
rect 20772 16204 20821 16232
rect 20772 16192 20778 16204
rect 20809 16201 20821 16204
rect 20855 16201 20867 16235
rect 20809 16195 20867 16201
rect 4157 16167 4215 16173
rect 4157 16133 4169 16167
rect 4203 16164 4215 16167
rect 5074 16164 5080 16176
rect 4203 16136 5080 16164
rect 4203 16133 4215 16136
rect 4157 16127 4215 16133
rect 5074 16124 5080 16136
rect 5132 16124 5138 16176
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 900 16068 1409 16096
rect 900 16056 906 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 3234 16056 3240 16108
rect 3292 16096 3298 16108
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 3292 16068 3985 16096
rect 3292 16056 3298 16068
rect 3973 16065 3985 16068
rect 4019 16065 4031 16099
rect 3973 16059 4031 16065
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16096 4859 16099
rect 5442 16096 5448 16108
rect 4847 16068 5448 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 6822 16056 6828 16108
rect 6880 16096 6886 16108
rect 7009 16099 7067 16105
rect 7009 16096 7021 16099
rect 6880 16068 7021 16096
rect 6880 16056 6886 16068
rect 7009 16065 7021 16068
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16096 7251 16099
rect 7282 16096 7288 16108
rect 7239 16068 7288 16096
rect 7239 16065 7251 16068
rect 7193 16059 7251 16065
rect 4246 15988 4252 16040
rect 4304 16028 4310 16040
rect 4709 16031 4767 16037
rect 4709 16028 4721 16031
rect 4304 16000 4721 16028
rect 4304 15988 4310 16000
rect 4709 15997 4721 16000
rect 4755 15997 4767 16031
rect 4709 15991 4767 15997
rect 5166 15988 5172 16040
rect 5224 15988 5230 16040
rect 7024 16028 7052 16059
rect 7282 16056 7288 16068
rect 7340 16096 7346 16108
rect 7653 16099 7711 16105
rect 7653 16096 7665 16099
rect 7340 16068 7665 16096
rect 7340 16056 7346 16068
rect 7653 16065 7665 16068
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 10042 16056 10048 16108
rect 10100 16056 10106 16108
rect 14090 16056 14096 16108
rect 14148 16056 14154 16108
rect 18506 16056 18512 16108
rect 18564 16056 18570 16108
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16096 20775 16099
rect 20763 16068 21864 16096
rect 20763 16065 20775 16068
rect 20717 16059 20775 16065
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7024 16000 7481 16028
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 7469 15991 7527 15997
rect 10321 16031 10379 16037
rect 10321 15997 10333 16031
rect 10367 16028 10379 16031
rect 11054 16028 11060 16040
rect 10367 16000 11060 16028
rect 10367 15997 10379 16000
rect 10321 15991 10379 15997
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 13722 16028 13728 16040
rect 13044 16000 13728 16028
rect 13044 15988 13050 16000
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18138 16028 18144 16040
rect 18012 16000 18144 16028
rect 18012 15988 18018 16000
rect 18138 15988 18144 16000
rect 18196 16028 18202 16040
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 18196 16000 18705 16028
rect 18196 15988 18202 16000
rect 18693 15997 18705 16000
rect 18739 16028 18751 16031
rect 19058 16028 19064 16040
rect 18739 16000 19064 16028
rect 18739 15997 18751 16000
rect 18693 15991 18751 15997
rect 19058 15988 19064 16000
rect 19116 16028 19122 16040
rect 20901 16031 20959 16037
rect 20901 16028 20913 16031
rect 19116 16000 20913 16028
rect 19116 15988 19122 16000
rect 20901 15997 20913 16000
rect 20947 16028 20959 16031
rect 21542 16028 21548 16040
rect 20947 16000 21548 16028
rect 20947 15997 20959 16000
rect 20901 15991 20959 15997
rect 21542 15988 21548 16000
rect 21600 15988 21606 16040
rect 21836 16037 21864 16068
rect 22186 16056 22192 16108
rect 22244 16056 22250 16108
rect 23658 16056 23664 16108
rect 23716 16056 23722 16108
rect 21821 16031 21879 16037
rect 21821 15997 21833 16031
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 22002 15988 22008 16040
rect 22060 16028 22066 16040
rect 22097 16031 22155 16037
rect 22097 16028 22109 16031
rect 22060 16000 22109 16028
rect 22060 15988 22066 16000
rect 22097 15997 22109 16000
rect 22143 15997 22155 16031
rect 22097 15991 22155 15997
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 7374 15960 7380 15972
rect 1627 15932 7380 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 7374 15920 7380 15932
rect 7432 15920 7438 15972
rect 6454 15852 6460 15904
rect 6512 15892 6518 15904
rect 7837 15895 7895 15901
rect 7837 15892 7849 15895
rect 6512 15864 7849 15892
rect 6512 15852 6518 15864
rect 7837 15861 7849 15864
rect 7883 15861 7895 15895
rect 7837 15855 7895 15861
rect 23477 15895 23535 15901
rect 23477 15861 23489 15895
rect 23523 15892 23535 15895
rect 23566 15892 23572 15904
rect 23523 15864 23572 15892
rect 23523 15861 23535 15864
rect 23477 15855 23535 15861
rect 23566 15852 23572 15864
rect 23624 15852 23630 15904
rect 1104 15802 24012 15824
rect 1104 15750 3813 15802
rect 3865 15750 3877 15802
rect 3929 15750 3941 15802
rect 3993 15750 4005 15802
rect 4057 15750 4069 15802
rect 4121 15750 9540 15802
rect 9592 15750 9604 15802
rect 9656 15750 9668 15802
rect 9720 15750 9732 15802
rect 9784 15750 9796 15802
rect 9848 15750 15267 15802
rect 15319 15750 15331 15802
rect 15383 15750 15395 15802
rect 15447 15750 15459 15802
rect 15511 15750 15523 15802
rect 15575 15750 20994 15802
rect 21046 15750 21058 15802
rect 21110 15750 21122 15802
rect 21174 15750 21186 15802
rect 21238 15750 21250 15802
rect 21302 15750 24012 15802
rect 1104 15728 24012 15750
rect 3234 15648 3240 15700
rect 3292 15648 3298 15700
rect 4982 15648 4988 15700
rect 5040 15648 5046 15700
rect 5074 15648 5080 15700
rect 5132 15648 5138 15700
rect 5368 15660 6868 15688
rect 1581 15623 1639 15629
rect 1581 15589 1593 15623
rect 1627 15620 1639 15623
rect 5368 15620 5396 15660
rect 1627 15592 5396 15620
rect 1627 15589 1639 15592
rect 1581 15583 1639 15589
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 6089 15623 6147 15629
rect 6089 15620 6101 15623
rect 5500 15592 6101 15620
rect 5500 15580 5506 15592
rect 6089 15589 6101 15592
rect 6135 15589 6147 15623
rect 6840 15620 6868 15660
rect 6914 15648 6920 15700
rect 6972 15648 6978 15700
rect 7745 15691 7803 15697
rect 7745 15657 7757 15691
rect 7791 15688 7803 15691
rect 8018 15688 8024 15700
rect 7791 15660 8024 15688
rect 7791 15657 7803 15660
rect 7745 15651 7803 15657
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 9858 15648 9864 15700
rect 9916 15688 9922 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 9916 15660 10057 15688
rect 9916 15648 9922 15660
rect 10045 15657 10057 15660
rect 10091 15657 10103 15691
rect 10045 15651 10103 15657
rect 14090 15648 14096 15700
rect 14148 15648 14154 15700
rect 19886 15648 19892 15700
rect 19944 15688 19950 15700
rect 20993 15691 21051 15697
rect 20993 15688 21005 15691
rect 19944 15660 21005 15688
rect 19944 15648 19950 15660
rect 20993 15657 21005 15660
rect 21039 15657 21051 15691
rect 20993 15651 21051 15657
rect 7006 15620 7012 15632
rect 6840 15592 7012 15620
rect 6089 15583 6147 15589
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 22186 15580 22192 15632
rect 22244 15580 22250 15632
rect 3605 15555 3663 15561
rect 3605 15521 3617 15555
rect 3651 15521 3663 15555
rect 3605 15515 3663 15521
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 5350 15552 5356 15564
rect 4479 15524 5356 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 3418 15444 3424 15496
rect 3476 15444 3482 15496
rect 3620 15428 3648 15515
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15552 6607 15555
rect 6638 15552 6644 15564
rect 6595 15524 6644 15552
rect 6595 15521 6607 15524
rect 6549 15515 6607 15521
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15552 6791 15555
rect 7282 15552 7288 15564
rect 6779 15524 7288 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15552 7619 15555
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7607 15524 8033 15552
rect 7607 15521 7619 15524
rect 7561 15515 7619 15521
rect 8021 15521 8033 15524
rect 8067 15552 8079 15555
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 8067 15524 8585 15552
rect 8067 15521 8079 15524
rect 8021 15515 8079 15521
rect 8573 15521 8585 15524
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 8754 15512 8760 15564
rect 8812 15512 8818 15564
rect 10689 15555 10747 15561
rect 10689 15521 10701 15555
rect 10735 15552 10747 15555
rect 11054 15552 11060 15564
rect 10735 15524 11060 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 14737 15555 14795 15561
rect 14737 15521 14749 15555
rect 14783 15552 14795 15555
rect 14826 15552 14832 15564
rect 14783 15524 14832 15552
rect 14783 15521 14795 15524
rect 14737 15515 14795 15521
rect 14826 15512 14832 15524
rect 14884 15512 14890 15564
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15552 15623 15555
rect 15654 15552 15660 15564
rect 15611 15524 15660 15552
rect 15611 15521 15623 15524
rect 15565 15515 15623 15521
rect 15654 15512 15660 15524
rect 15712 15512 15718 15564
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18874 15552 18880 15564
rect 18187 15524 18880 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18874 15512 18880 15524
rect 18932 15512 18938 15564
rect 21542 15512 21548 15564
rect 21600 15512 21606 15564
rect 4246 15444 4252 15496
rect 4304 15484 4310 15496
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 4304 15456 5273 15484
rect 4304 15444 4310 15456
rect 5261 15453 5273 15456
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 6319 15456 6684 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 3602 15376 3608 15428
rect 3660 15416 3666 15428
rect 3789 15419 3847 15425
rect 3789 15416 3801 15419
rect 3660 15388 3801 15416
rect 3660 15376 3666 15388
rect 3789 15385 3801 15388
rect 3835 15385 3847 15419
rect 3973 15419 4031 15425
rect 3973 15416 3985 15419
rect 3789 15379 3847 15385
rect 3896 15388 3985 15416
rect 3418 15308 3424 15360
rect 3476 15348 3482 15360
rect 3896 15348 3924 15388
rect 3973 15385 3985 15388
rect 4019 15385 4031 15419
rect 3973 15379 4031 15385
rect 6454 15376 6460 15428
rect 6512 15376 6518 15428
rect 6656 15416 6684 15456
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 7193 15487 7251 15493
rect 7193 15484 7205 15487
rect 6880 15456 7205 15484
rect 6880 15444 6886 15456
rect 7193 15453 7205 15456
rect 7239 15453 7251 15487
rect 7193 15447 7251 15453
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 8772 15484 8800 15512
rect 8159 15456 8800 15484
rect 15381 15487 15439 15493
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 15381 15453 15393 15487
rect 15427 15484 15439 15487
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 15427 15456 15761 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 15749 15453 15761 15456
rect 15795 15453 15807 15487
rect 15749 15447 15807 15453
rect 17954 15444 17960 15496
rect 18012 15444 18018 15496
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 23382 15444 23388 15496
rect 23440 15484 23446 15496
rect 23661 15487 23719 15493
rect 23661 15484 23673 15487
rect 23440 15456 23673 15484
rect 23440 15444 23446 15456
rect 23661 15453 23673 15456
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 8389 15419 8447 15425
rect 8389 15416 8401 15419
rect 6656 15388 8401 15416
rect 8389 15385 8401 15388
rect 8435 15385 8447 15419
rect 8389 15379 8447 15385
rect 10413 15419 10471 15425
rect 10413 15385 10425 15419
rect 10459 15416 10471 15419
rect 10686 15416 10692 15428
rect 10459 15388 10692 15416
rect 10459 15385 10471 15388
rect 10413 15379 10471 15385
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 3476 15320 3924 15348
rect 4157 15351 4215 15357
rect 3476 15308 3482 15320
rect 4157 15317 4169 15351
rect 4203 15348 4215 15351
rect 4525 15351 4583 15357
rect 4525 15348 4537 15351
rect 4203 15320 4537 15348
rect 4203 15317 4215 15320
rect 4157 15311 4215 15317
rect 4525 15317 4537 15320
rect 4571 15317 4583 15351
rect 4525 15311 4583 15317
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15348 4675 15351
rect 4798 15348 4804 15360
rect 4663 15320 4804 15348
rect 4663 15317 4675 15320
rect 4617 15311 4675 15317
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 10505 15351 10563 15357
rect 10505 15317 10517 15351
rect 10551 15348 10563 15351
rect 10594 15348 10600 15360
rect 10551 15320 10600 15348
rect 10551 15317 10563 15320
rect 10505 15311 10563 15317
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 14458 15308 14464 15360
rect 14516 15308 14522 15360
rect 14553 15351 14611 15357
rect 14553 15317 14565 15351
rect 14599 15348 14611 15351
rect 14921 15351 14979 15357
rect 14921 15348 14933 15351
rect 14599 15320 14933 15348
rect 14599 15317 14611 15320
rect 14553 15311 14611 15317
rect 14921 15317 14933 15320
rect 14967 15317 14979 15351
rect 14921 15311 14979 15317
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15289 15351 15347 15357
rect 15289 15348 15301 15351
rect 15252 15320 15301 15348
rect 15252 15308 15258 15320
rect 15289 15317 15301 15320
rect 15335 15317 15347 15351
rect 15289 15311 15347 15317
rect 17126 15308 17132 15360
rect 17184 15348 17190 15360
rect 17773 15351 17831 15357
rect 17773 15348 17785 15351
rect 17184 15320 17785 15348
rect 17184 15308 17190 15320
rect 17773 15317 17785 15320
rect 17819 15317 17831 15351
rect 17773 15311 17831 15317
rect 21358 15308 21364 15360
rect 21416 15308 21422 15360
rect 21450 15308 21456 15360
rect 21508 15308 21514 15360
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 21821 15351 21879 15357
rect 21821 15348 21833 15351
rect 21600 15320 21833 15348
rect 21600 15308 21606 15320
rect 21821 15317 21833 15320
rect 21867 15317 21879 15351
rect 21821 15311 21879 15317
rect 23477 15351 23535 15357
rect 23477 15317 23489 15351
rect 23523 15348 23535 15351
rect 23658 15348 23664 15360
rect 23523 15320 23664 15348
rect 23523 15317 23535 15320
rect 23477 15311 23535 15317
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 1104 15258 24012 15280
rect 1104 15206 4473 15258
rect 4525 15206 4537 15258
rect 4589 15206 4601 15258
rect 4653 15206 4665 15258
rect 4717 15206 4729 15258
rect 4781 15206 10200 15258
rect 10252 15206 10264 15258
rect 10316 15206 10328 15258
rect 10380 15206 10392 15258
rect 10444 15206 10456 15258
rect 10508 15206 15927 15258
rect 15979 15206 15991 15258
rect 16043 15206 16055 15258
rect 16107 15206 16119 15258
rect 16171 15206 16183 15258
rect 16235 15206 21654 15258
rect 21706 15206 21718 15258
rect 21770 15206 21782 15258
rect 21834 15206 21846 15258
rect 21898 15206 21910 15258
rect 21962 15206 24012 15258
rect 1104 15184 24012 15206
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4798 15144 4804 15156
rect 4755 15116 4804 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 7009 15147 7067 15153
rect 7009 15113 7021 15147
rect 7055 15144 7067 15147
rect 7282 15144 7288 15156
rect 7055 15116 7288 15144
rect 7055 15113 7067 15116
rect 7009 15107 7067 15113
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 7374 15104 7380 15156
rect 7432 15104 7438 15156
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 9309 15147 9367 15153
rect 9309 15144 9321 15147
rect 8812 15116 9321 15144
rect 8812 15104 8818 15116
rect 9309 15113 9321 15116
rect 9355 15113 9367 15147
rect 9309 15107 9367 15113
rect 10594 15104 10600 15156
rect 10652 15104 10658 15156
rect 10686 15104 10692 15156
rect 10744 15104 10750 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18417 15147 18475 15153
rect 18417 15144 18429 15147
rect 18104 15116 18429 15144
rect 18104 15104 18110 15116
rect 18417 15113 18429 15116
rect 18463 15113 18475 15147
rect 18417 15107 18475 15113
rect 20809 15147 20867 15153
rect 20809 15113 20821 15147
rect 20855 15144 20867 15147
rect 21358 15144 21364 15156
rect 20855 15116 21364 15144
rect 20855 15113 20867 15116
rect 20809 15107 20867 15113
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 8662 15076 8668 15088
rect 7668 15048 8668 15076
rect 3602 14968 3608 15020
rect 3660 15008 3666 15020
rect 3881 15011 3939 15017
rect 3881 15008 3893 15011
rect 3660 14980 3893 15008
rect 3660 14968 3666 14980
rect 3881 14977 3893 14980
rect 3927 15008 3939 15011
rect 3927 14980 4384 15008
rect 3927 14977 3939 14980
rect 3881 14971 3939 14977
rect 3418 14900 3424 14952
rect 3476 14940 3482 14952
rect 3694 14940 3700 14952
rect 3476 14912 3700 14940
rect 3476 14900 3482 14912
rect 3694 14900 3700 14912
rect 3752 14940 3758 14952
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 3752 14912 3801 14940
rect 3752 14900 3758 14912
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 3804 14872 3832 14903
rect 4246 14900 4252 14952
rect 4304 14900 4310 14952
rect 4356 14949 4384 14980
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 7668 15008 7696 15048
rect 8662 15036 8668 15048
rect 8720 15076 8726 15088
rect 12434 15076 12440 15088
rect 8720 15048 12440 15076
rect 8720 15036 8726 15048
rect 12434 15036 12440 15048
rect 12492 15076 12498 15088
rect 13078 15076 13084 15088
rect 12492 15048 13084 15076
rect 12492 15036 12498 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 21453 15079 21511 15085
rect 18012 15048 18828 15076
rect 18012 15036 18018 15048
rect 5316 14980 7696 15008
rect 5316 14968 5322 14980
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 4540 14872 4568 14903
rect 7466 14900 7472 14952
rect 7524 14900 7530 14952
rect 7668 14949 7696 14980
rect 9398 14968 9404 15020
rect 9456 15008 9462 15020
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9456 14980 9505 15008
rect 9456 14968 9462 14980
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 15008 9735 15011
rect 9769 15011 9827 15017
rect 9769 15008 9781 15011
rect 9723 14980 9781 15008
rect 9723 14977 9735 14980
rect 9677 14971 9735 14977
rect 9769 14977 9781 14980
rect 9815 14977 9827 15011
rect 10229 15011 10287 15017
rect 10229 15008 10241 15011
rect 9769 14971 9827 14977
rect 10152 14980 10241 15008
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 3804 14844 4568 14872
rect 9968 14804 9996 14903
rect 10152 14881 10180 14980
rect 10229 14977 10241 14980
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 10428 14940 10456 14971
rect 11882 14968 11888 15020
rect 11940 15017 11946 15020
rect 11940 15011 11978 15017
rect 11966 14977 11978 15011
rect 11940 14971 11978 14977
rect 11940 14968 11946 14971
rect 15654 14968 15660 15020
rect 15712 15008 15718 15020
rect 17862 15008 17868 15020
rect 15712 14980 17868 15008
rect 15712 14968 15718 14980
rect 10870 14940 10876 14952
rect 10428 14912 10876 14940
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 17788 14949 17816 14980
rect 17862 14968 17868 14980
rect 17920 14968 17926 15020
rect 18046 14968 18052 15020
rect 18104 14968 18110 15020
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14940 17371 14943
rect 17773 14943 17831 14949
rect 17359 14912 17724 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 10137 14875 10195 14881
rect 10137 14841 10149 14875
rect 10183 14872 10195 14875
rect 10226 14872 10232 14884
rect 10183 14844 10232 14872
rect 10183 14841 10195 14844
rect 10137 14835 10195 14841
rect 10226 14832 10232 14844
rect 10284 14872 10290 14884
rect 11057 14875 11115 14881
rect 11057 14872 11069 14875
rect 10284 14844 11069 14872
rect 10284 14832 10290 14844
rect 11057 14841 11069 14844
rect 11103 14872 11115 14875
rect 12342 14872 12348 14884
rect 11103 14844 12348 14872
rect 11103 14841 11115 14844
rect 11057 14835 11115 14841
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 17497 14875 17555 14881
rect 17497 14841 17509 14875
rect 17543 14872 17555 14875
rect 17586 14872 17592 14884
rect 17543 14844 17592 14872
rect 17543 14841 17555 14844
rect 17497 14835 17555 14841
rect 17586 14832 17592 14844
rect 17644 14832 17650 14884
rect 17696 14872 17724 14912
rect 17773 14909 17785 14943
rect 17819 14909 17831 14943
rect 17773 14903 17831 14909
rect 17957 14943 18015 14949
rect 17957 14909 17969 14943
rect 18003 14940 18015 14943
rect 18414 14940 18420 14952
rect 18003 14912 18420 14940
rect 18003 14909 18015 14912
rect 17957 14903 18015 14909
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 18506 14900 18512 14952
rect 18564 14900 18570 14952
rect 18800 14949 18828 15048
rect 21453 15045 21465 15079
rect 21499 15076 21511 15079
rect 21542 15076 21548 15088
rect 21499 15048 21548 15076
rect 21499 15045 21511 15048
rect 21453 15039 21511 15045
rect 21542 15036 21548 15048
rect 21600 15036 21606 15088
rect 22925 15079 22983 15085
rect 21744 15048 22140 15076
rect 18874 14968 18880 15020
rect 18932 15008 18938 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 18932 14980 21281 15008
rect 18932 14968 18938 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21634 14968 21640 15020
rect 21692 14968 21698 15020
rect 18785 14943 18843 14949
rect 18785 14909 18797 14943
rect 18831 14909 18843 14943
rect 18785 14903 18843 14909
rect 20993 14943 21051 14949
rect 20993 14909 21005 14943
rect 21039 14940 21051 14943
rect 21744 14940 21772 15048
rect 22112 14952 22140 15048
rect 22925 15045 22937 15079
rect 22971 15076 22983 15079
rect 22971 15048 23612 15076
rect 22971 15045 22983 15048
rect 22925 15039 22983 15045
rect 23584 15020 23612 15048
rect 23566 15017 23572 15020
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 23017 15011 23075 15017
rect 23017 14977 23029 15011
rect 23063 15008 23075 15011
rect 23431 15011 23489 15017
rect 23431 15008 23443 15011
rect 23063 14980 23443 15008
rect 23063 14977 23075 14980
rect 23017 14971 23075 14977
rect 23431 14977 23443 14980
rect 23477 14977 23489 15011
rect 23431 14971 23489 14977
rect 23534 15011 23572 15017
rect 23534 14977 23546 15011
rect 23534 14971 23572 14977
rect 21039 14912 21772 14940
rect 21821 14943 21879 14949
rect 21039 14909 21051 14912
rect 20993 14903 21051 14909
rect 21821 14909 21833 14943
rect 21867 14940 21879 14943
rect 22002 14940 22008 14952
rect 21867 14912 22008 14940
rect 21867 14909 21879 14912
rect 21821 14903 21879 14909
rect 22002 14900 22008 14912
rect 22060 14900 22066 14952
rect 22094 14900 22100 14952
rect 22152 14900 22158 14952
rect 17862 14872 17868 14884
rect 17696 14844 17868 14872
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 21177 14875 21235 14881
rect 21177 14841 21189 14875
rect 21223 14872 21235 14875
rect 22204 14872 22232 14971
rect 23566 14968 23572 14971
rect 23624 14968 23630 15020
rect 23201 14943 23259 14949
rect 23201 14909 23213 14943
rect 23247 14940 23259 14943
rect 23290 14940 23296 14952
rect 23247 14912 23296 14940
rect 23247 14909 23259 14912
rect 23201 14903 23259 14909
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 22557 14875 22615 14881
rect 22557 14872 22569 14875
rect 21223 14844 22094 14872
rect 21223 14841 21235 14844
rect 21177 14835 21235 14841
rect 10870 14804 10876 14816
rect 9968 14776 10876 14804
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 12023 14807 12081 14813
rect 12023 14773 12035 14807
rect 12069 14804 12081 14807
rect 12802 14804 12808 14816
rect 12069 14776 12808 14804
rect 12069 14773 12081 14776
rect 12023 14767 12081 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 17129 14807 17187 14813
rect 17129 14773 17141 14807
rect 17175 14804 17187 14807
rect 17310 14804 17316 14816
rect 17175 14776 17316 14804
rect 17175 14773 17187 14776
rect 17129 14767 17187 14773
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 22066 14804 22094 14844
rect 22204 14844 22569 14872
rect 22204 14804 22232 14844
rect 22557 14841 22569 14844
rect 22603 14841 22615 14875
rect 22557 14835 22615 14841
rect 22278 14804 22284 14816
rect 22066 14776 22284 14804
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 1104 14714 24012 14736
rect 1104 14662 3813 14714
rect 3865 14662 3877 14714
rect 3929 14662 3941 14714
rect 3993 14662 4005 14714
rect 4057 14662 4069 14714
rect 4121 14662 9540 14714
rect 9592 14662 9604 14714
rect 9656 14662 9668 14714
rect 9720 14662 9732 14714
rect 9784 14662 9796 14714
rect 9848 14662 15267 14714
rect 15319 14662 15331 14714
rect 15383 14662 15395 14714
rect 15447 14662 15459 14714
rect 15511 14662 15523 14714
rect 15575 14662 20994 14714
rect 21046 14662 21058 14714
rect 21110 14662 21122 14714
rect 21174 14662 21186 14714
rect 21238 14662 21250 14714
rect 21302 14662 24012 14714
rect 1104 14640 24012 14662
rect 3602 14560 3608 14612
rect 3660 14560 3666 14612
rect 3694 14560 3700 14612
rect 3752 14600 3758 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 3752 14572 4261 14600
rect 3752 14560 3758 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 6638 14560 6644 14612
rect 6696 14560 6702 14612
rect 7466 14560 7472 14612
rect 7524 14609 7530 14612
rect 7524 14603 7573 14609
rect 7524 14569 7527 14603
rect 7561 14569 7573 14603
rect 7524 14563 7573 14569
rect 7524 14560 7530 14563
rect 9398 14560 9404 14612
rect 9456 14560 9462 14612
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 10505 14603 10563 14609
rect 10505 14600 10517 14603
rect 10100 14572 10517 14600
rect 10100 14560 10106 14572
rect 10505 14569 10517 14572
rect 10551 14569 10563 14603
rect 10505 14563 10563 14569
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 10928 14572 11529 14600
rect 10928 14560 10934 14572
rect 11517 14569 11529 14572
rect 11563 14569 11575 14603
rect 11517 14563 11575 14569
rect 12342 14560 12348 14612
rect 12400 14560 12406 14612
rect 14458 14560 14464 14612
rect 14516 14600 14522 14612
rect 14829 14603 14887 14609
rect 14829 14600 14841 14603
rect 14516 14572 14841 14600
rect 14516 14560 14522 14572
rect 14829 14569 14841 14572
rect 14875 14569 14887 14603
rect 14829 14563 14887 14569
rect 15102 14560 15108 14612
rect 15160 14560 15166 14612
rect 17954 14560 17960 14612
rect 18012 14560 18018 14612
rect 18414 14560 18420 14612
rect 18472 14560 18478 14612
rect 21450 14560 21456 14612
rect 21508 14560 21514 14612
rect 21634 14560 21640 14612
rect 21692 14600 21698 14612
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 21692 14572 21925 14600
rect 21692 14560 21698 14572
rect 21913 14569 21925 14572
rect 21959 14569 21971 14603
rect 23658 14600 23664 14612
rect 21913 14563 21971 14569
rect 22066 14572 23664 14600
rect 9861 14535 9919 14541
rect 9861 14532 9873 14535
rect 3068 14504 7236 14532
rect 3068 14473 3096 14504
rect 7208 14476 7236 14504
rect 9600 14504 9873 14532
rect 3053 14467 3111 14473
rect 3053 14433 3065 14467
rect 3099 14433 3111 14467
rect 3053 14427 3111 14433
rect 4893 14467 4951 14473
rect 4893 14433 4905 14467
rect 4939 14464 4951 14467
rect 5074 14464 5080 14476
rect 4939 14436 5080 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 7190 14424 7196 14476
rect 7248 14424 7254 14476
rect 9600 14473 9628 14504
rect 9861 14501 9873 14504
rect 9907 14532 9919 14535
rect 9907 14504 10824 14532
rect 9907 14501 9919 14504
rect 9861 14495 9919 14501
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14464 9827 14467
rect 9950 14464 9956 14476
rect 9815 14436 9956 14464
rect 9815 14433 9827 14436
rect 9769 14427 9827 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14464 10379 14467
rect 10686 14464 10692 14476
rect 10367 14436 10692 14464
rect 10367 14433 10379 14436
rect 10321 14427 10379 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 10796 14473 10824 14504
rect 11054 14492 11060 14544
rect 11112 14532 11118 14544
rect 15654 14532 15660 14544
rect 11112 14504 15660 14532
rect 11112 14492 11118 14504
rect 10781 14467 10839 14473
rect 10781 14433 10793 14467
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 12161 14467 12219 14473
rect 12161 14433 12173 14467
rect 12207 14464 12219 14467
rect 12434 14464 12440 14476
rect 12207 14436 12440 14464
rect 12207 14433 12219 14436
rect 12161 14427 12219 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 12802 14424 12808 14476
rect 12860 14424 12866 14476
rect 12986 14424 12992 14476
rect 13044 14424 13050 14476
rect 14200 14473 14228 14504
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 22066 14532 22094 14572
rect 23658 14560 23664 14572
rect 23716 14560 23722 14612
rect 19628 14504 22094 14532
rect 14185 14467 14243 14473
rect 14185 14433 14197 14467
rect 14231 14433 14243 14467
rect 14185 14427 14243 14433
rect 15562 14424 15568 14476
rect 15620 14424 15626 14476
rect 17681 14467 17739 14473
rect 17681 14433 17693 14467
rect 17727 14464 17739 14467
rect 17727 14436 18276 14464
rect 17727 14433 17739 14436
rect 17681 14427 17739 14433
rect 842 14356 848 14408
rect 900 14396 906 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 900 14368 1409 14396
rect 900 14356 906 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 3237 14399 3295 14405
rect 3237 14396 3249 14399
rect 1397 14359 1455 14365
rect 2746 14368 3249 14396
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 2746 14260 2774 14368
rect 3237 14365 3249 14368
rect 3283 14396 3295 14399
rect 3922 14399 3980 14405
rect 3922 14396 3934 14399
rect 3283 14368 3934 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3922 14365 3934 14368
rect 3968 14365 3980 14399
rect 5194 14399 5252 14405
rect 5194 14396 5206 14399
rect 3922 14359 3980 14365
rect 4632 14368 5206 14396
rect 3145 14331 3203 14337
rect 3145 14297 3157 14331
rect 3191 14328 3203 14331
rect 3835 14331 3893 14337
rect 3835 14328 3847 14331
rect 3191 14300 3847 14328
rect 3191 14297 3203 14300
rect 3145 14291 3203 14297
rect 3835 14297 3847 14300
rect 3881 14297 3893 14331
rect 3835 14291 3893 14297
rect 1627 14232 2774 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 4632 14269 4660 14368
rect 5194 14365 5206 14368
rect 5240 14365 5252 14399
rect 5194 14359 5252 14365
rect 7006 14356 7012 14408
rect 7064 14356 7070 14408
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7586 14399 7644 14405
rect 7586 14396 7598 14399
rect 7432 14368 7598 14396
rect 7432 14356 7438 14368
rect 7586 14365 7598 14368
rect 7632 14365 7644 14399
rect 7862 14399 7920 14405
rect 7862 14396 7874 14399
rect 7586 14359 7644 14365
rect 7760 14368 7874 14396
rect 7024 14328 7052 14356
rect 7760 14328 7788 14368
rect 7862 14365 7874 14368
rect 7908 14365 7920 14399
rect 7862 14359 7920 14365
rect 10226 14356 10232 14408
rect 10284 14356 10290 14408
rect 10873 14399 10931 14405
rect 10873 14365 10885 14399
rect 10919 14365 10931 14399
rect 10873 14359 10931 14365
rect 7024 14300 7788 14328
rect 9950 14288 9956 14340
rect 10008 14328 10014 14340
rect 10888 14328 10916 14359
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 13541 14399 13599 14405
rect 11940 14368 12434 14396
rect 11940 14356 11946 14368
rect 10008 14300 10916 14328
rect 12406 14328 12434 14368
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13814 14396 13820 14408
rect 13587 14368 13820 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 15654 14396 15660 14408
rect 15519 14368 15660 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15654 14356 15660 14368
rect 15712 14396 15718 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 15712 14368 16957 14396
rect 15712 14356 15718 14368
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 17126 14356 17132 14408
rect 17184 14356 17190 14408
rect 17310 14356 17316 14408
rect 17368 14356 17374 14408
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 18049 14399 18107 14405
rect 18049 14396 18061 14399
rect 17644 14368 18061 14396
rect 17644 14356 17650 14368
rect 18049 14365 18061 14368
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 12713 14331 12771 14337
rect 12713 14328 12725 14331
rect 12406 14300 12725 14328
rect 10008 14288 10014 14300
rect 12713 14297 12725 14300
rect 12759 14297 12771 14331
rect 12713 14291 12771 14297
rect 13725 14331 13783 14337
rect 13725 14297 13737 14331
rect 13771 14328 13783 14331
rect 14090 14328 14096 14340
rect 13771 14300 14096 14328
rect 13771 14297 13783 14300
rect 13725 14291 13783 14297
rect 14090 14288 14096 14300
rect 14148 14288 14154 14340
rect 18248 14337 18276 14436
rect 19628 14405 19656 14504
rect 22278 14492 22284 14544
rect 22336 14492 22342 14544
rect 19889 14467 19947 14473
rect 19889 14433 19901 14467
rect 19935 14433 19947 14467
rect 22296 14464 22324 14492
rect 23106 14464 23112 14476
rect 19889 14427 19947 14433
rect 21560 14436 22324 14464
rect 22388 14436 23112 14464
rect 18928 14399 18986 14405
rect 18928 14365 18940 14399
rect 18974 14396 18986 14399
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 18974 14368 19625 14396
rect 18974 14365 18986 14368
rect 18928 14359 18986 14365
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 18233 14331 18291 14337
rect 18233 14297 18245 14331
rect 18279 14297 18291 14331
rect 18233 14291 18291 14297
rect 19015 14331 19073 14337
rect 19015 14297 19027 14331
rect 19061 14328 19073 14331
rect 19705 14331 19763 14337
rect 19705 14328 19717 14331
rect 19061 14300 19717 14328
rect 19061 14297 19073 14300
rect 19015 14291 19073 14297
rect 19705 14297 19717 14300
rect 19751 14297 19763 14331
rect 19705 14291 19763 14297
rect 4617 14263 4675 14269
rect 4617 14260 4629 14263
rect 4396 14232 4629 14260
rect 4396 14220 4402 14232
rect 4617 14229 4629 14232
rect 4663 14229 4675 14263
rect 4617 14223 4675 14229
rect 4709 14263 4767 14269
rect 4709 14229 4721 14263
rect 4755 14260 4767 14263
rect 5123 14263 5181 14269
rect 5123 14260 5135 14263
rect 4755 14232 5135 14260
rect 4755 14229 4767 14232
rect 4709 14223 4767 14229
rect 5123 14229 5135 14232
rect 5169 14229 5181 14263
rect 5123 14223 5181 14229
rect 7101 14263 7159 14269
rect 7101 14229 7113 14263
rect 7147 14260 7159 14263
rect 7791 14263 7849 14269
rect 7791 14260 7803 14263
rect 7147 14232 7803 14260
rect 7147 14229 7159 14232
rect 7101 14223 7159 14229
rect 7791 14229 7803 14232
rect 7837 14229 7849 14263
rect 7791 14223 7849 14229
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 11885 14263 11943 14269
rect 11885 14260 11897 14263
rect 11848 14232 11897 14260
rect 11848 14220 11854 14232
rect 11885 14229 11897 14232
rect 11931 14229 11943 14263
rect 11885 14223 11943 14229
rect 11974 14220 11980 14272
rect 12032 14220 12038 14272
rect 13909 14263 13967 14269
rect 13909 14229 13921 14263
rect 13955 14260 13967 14263
rect 14369 14263 14427 14269
rect 14369 14260 14381 14263
rect 13955 14232 14381 14260
rect 13955 14229 13967 14232
rect 13909 14223 13967 14229
rect 14369 14229 14381 14232
rect 14415 14229 14427 14263
rect 14369 14223 14427 14229
rect 14458 14220 14464 14272
rect 14516 14220 14522 14272
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 18248 14260 18276 14291
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 17920 14232 19257 14260
rect 17920 14220 17926 14232
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 19904 14260 19932 14427
rect 21560 14328 21588 14436
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14396 21695 14399
rect 21683 14368 21956 14396
rect 21683 14365 21695 14368
rect 21637 14359 21695 14365
rect 21821 14331 21879 14337
rect 21821 14328 21833 14331
rect 21560 14300 21833 14328
rect 21821 14297 21833 14300
rect 21867 14297 21879 14331
rect 21928 14328 21956 14368
rect 22094 14356 22100 14408
rect 22152 14356 22158 14408
rect 22186 14356 22192 14408
rect 22244 14396 22250 14408
rect 22388 14396 22416 14436
rect 23106 14424 23112 14436
rect 23164 14424 23170 14476
rect 22244 14368 22416 14396
rect 22925 14399 22983 14405
rect 22244 14356 22250 14368
rect 22925 14365 22937 14399
rect 22971 14396 22983 14399
rect 23474 14396 23480 14408
rect 23532 14405 23538 14408
rect 23532 14399 23560 14405
rect 22971 14368 23480 14396
rect 22971 14365 22983 14368
rect 22925 14359 22983 14365
rect 23474 14356 23480 14368
rect 23548 14365 23560 14399
rect 23532 14359 23560 14365
rect 23532 14356 23538 14359
rect 22112 14328 22140 14356
rect 21928 14300 22600 14328
rect 21821 14291 21879 14297
rect 22186 14260 22192 14272
rect 19904 14232 22192 14260
rect 19245 14223 19303 14229
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 22572 14269 22600 14300
rect 22557 14263 22615 14269
rect 22557 14229 22569 14263
rect 22603 14229 22615 14263
rect 22557 14223 22615 14229
rect 23017 14263 23075 14269
rect 23017 14229 23029 14263
rect 23063 14260 23075 14263
rect 23431 14263 23489 14269
rect 23431 14260 23443 14263
rect 23063 14232 23443 14260
rect 23063 14229 23075 14232
rect 23017 14223 23075 14229
rect 23431 14229 23443 14232
rect 23477 14229 23489 14263
rect 23431 14223 23489 14229
rect 1104 14170 24012 14192
rect 1104 14118 4473 14170
rect 4525 14118 4537 14170
rect 4589 14118 4601 14170
rect 4653 14118 4665 14170
rect 4717 14118 4729 14170
rect 4781 14118 10200 14170
rect 10252 14118 10264 14170
rect 10316 14118 10328 14170
rect 10380 14118 10392 14170
rect 10444 14118 10456 14170
rect 10508 14118 15927 14170
rect 15979 14118 15991 14170
rect 16043 14118 16055 14170
rect 16107 14118 16119 14170
rect 16171 14118 16183 14170
rect 16235 14118 21654 14170
rect 21706 14118 21718 14170
rect 21770 14118 21782 14170
rect 21834 14118 21846 14170
rect 21898 14118 21910 14170
rect 21962 14118 24012 14170
rect 1104 14096 24012 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 4338 14056 4344 14068
rect 1627 14028 4344 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 11974 14065 11980 14068
rect 11931 14059 11980 14065
rect 11931 14025 11943 14059
rect 11977 14025 11980 14059
rect 11931 14019 11980 14025
rect 11974 14016 11980 14019
rect 12032 14016 12038 14068
rect 14185 14059 14243 14065
rect 14185 14025 14197 14059
rect 14231 14056 14243 14059
rect 14458 14056 14464 14068
rect 14231 14028 14464 14056
rect 14231 14025 14243 14028
rect 14185 14019 14243 14025
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 17586 14016 17592 14068
rect 17644 14016 17650 14068
rect 18046 14016 18052 14068
rect 18104 14016 18110 14068
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 12002 13923 12060 13929
rect 12002 13920 12014 13923
rect 11848 13892 12014 13920
rect 11848 13880 11854 13892
rect 12002 13889 12014 13892
rect 12048 13889 12060 13923
rect 14461 13923 14519 13929
rect 14461 13920 14473 13923
rect 12002 13883 12060 13889
rect 13832 13892 14473 13920
rect 13832 13864 13860 13892
rect 14461 13889 14473 13892
rect 14507 13889 14519 13923
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 14461 13883 14519 13889
rect 14844 13892 15485 13920
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14090 13852 14096 13864
rect 14047 13824 14096 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14090 13812 14096 13824
rect 14148 13852 14154 13864
rect 14844 13861 14872 13892
rect 15473 13889 15485 13892
rect 15519 13920 15531 13923
rect 15562 13920 15568 13932
rect 15519 13892 15568 13920
rect 15519 13889 15531 13892
rect 15473 13883 15531 13889
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 14369 13855 14427 13861
rect 14369 13852 14381 13855
rect 14148 13824 14381 13852
rect 14148 13812 14154 13824
rect 14369 13821 14381 13824
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13821 14887 13855
rect 14829 13815 14887 13821
rect 15654 13812 15660 13864
rect 15712 13812 15718 13864
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13821 17095 13855
rect 17037 13815 17095 13821
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 12986 13784 12992 13796
rect 7248 13756 12992 13784
rect 7248 13744 7254 13756
rect 12986 13744 12992 13756
rect 13044 13744 13050 13796
rect 17052 13728 17080 13815
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 17236 13796 17264 13883
rect 17604 13852 17632 14016
rect 17862 13880 17868 13932
rect 17920 13880 17926 13932
rect 23382 13880 23388 13932
rect 23440 13880 23446 13932
rect 23658 13880 23664 13932
rect 23716 13880 23722 13932
rect 17681 13855 17739 13861
rect 17681 13852 17693 13855
rect 17604 13824 17693 13852
rect 17681 13821 17693 13824
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 17972 13824 23520 13852
rect 17218 13744 17224 13796
rect 17276 13784 17282 13796
rect 17972 13784 18000 13824
rect 23492 13793 23520 13824
rect 17276 13756 18000 13784
rect 23477 13787 23535 13793
rect 17276 13744 17282 13756
rect 23477 13753 23489 13787
rect 23523 13753 23535 13787
rect 23477 13747 23535 13753
rect 15289 13719 15347 13725
rect 15289 13685 15301 13719
rect 15335 13716 15347 13719
rect 15746 13716 15752 13728
rect 15335 13688 15752 13716
rect 15335 13685 15347 13688
rect 15289 13679 15347 13685
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 17034 13676 17040 13728
rect 17092 13676 17098 13728
rect 23198 13676 23204 13728
rect 23256 13676 23262 13728
rect 1104 13626 24012 13648
rect 1104 13574 3813 13626
rect 3865 13574 3877 13626
rect 3929 13574 3941 13626
rect 3993 13574 4005 13626
rect 4057 13574 4069 13626
rect 4121 13574 9540 13626
rect 9592 13574 9604 13626
rect 9656 13574 9668 13626
rect 9720 13574 9732 13626
rect 9784 13574 9796 13626
rect 9848 13574 15267 13626
rect 15319 13574 15331 13626
rect 15383 13574 15395 13626
rect 15447 13574 15459 13626
rect 15511 13574 15523 13626
rect 15575 13574 20994 13626
rect 21046 13574 21058 13626
rect 21110 13574 21122 13626
rect 21174 13574 21186 13626
rect 21238 13574 21250 13626
rect 21302 13574 24012 13626
rect 1104 13552 24012 13574
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 13872 13484 14412 13512
rect 13872 13472 13878 13484
rect 14384 13453 14412 13484
rect 17126 13472 17132 13524
rect 17184 13521 17190 13524
rect 17184 13515 17233 13521
rect 17184 13481 17187 13515
rect 17221 13481 17233 13515
rect 17184 13475 17233 13481
rect 17184 13472 17190 13475
rect 14369 13447 14427 13453
rect 14369 13413 14381 13447
rect 14415 13413 14427 13447
rect 23198 13444 23204 13456
rect 14369 13407 14427 13413
rect 15396 13416 23204 13444
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13173 13379 13231 13385
rect 13173 13376 13185 13379
rect 13044 13348 13185 13376
rect 13044 13336 13050 13348
rect 13173 13345 13185 13348
rect 13219 13376 13231 13379
rect 13262 13376 13268 13388
rect 13219 13348 13268 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 14553 13379 14611 13385
rect 14553 13376 14565 13379
rect 14148 13348 14565 13376
rect 14148 13336 14154 13348
rect 14553 13345 14565 13348
rect 14599 13345 14611 13379
rect 14553 13339 14611 13345
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 7006 13317 7012 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 900 13280 1409 13308
rect 900 13268 906 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 6984 13311 7012 13317
rect 6984 13277 6996 13311
rect 6984 13271 7012 13277
rect 7006 13268 7012 13271
rect 7064 13268 7070 13320
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13308 13507 13311
rect 14242 13311 14300 13317
rect 14242 13308 14254 13311
rect 13495 13280 14254 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 14242 13277 14254 13280
rect 14288 13308 14300 13311
rect 15396 13308 15424 13416
rect 23198 13404 23204 13416
rect 23256 13404 23262 13456
rect 23477 13447 23535 13453
rect 23477 13413 23489 13447
rect 23523 13413 23535 13447
rect 23477 13407 23535 13413
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13376 19671 13379
rect 19978 13376 19984 13388
rect 19659 13348 19984 13376
rect 19659 13345 19671 13348
rect 19613 13339 19671 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 14288 13280 15424 13308
rect 15473 13311 15531 13317
rect 14288 13277 14300 13280
rect 14242 13271 14300 13277
rect 15473 13277 15485 13311
rect 15519 13308 15531 13311
rect 15746 13308 15752 13320
rect 15519 13280 15752 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 17218 13268 17224 13320
rect 17276 13317 17282 13320
rect 17276 13311 17304 13317
rect 17292 13277 17304 13311
rect 17276 13271 17304 13277
rect 17276 13268 17282 13271
rect 19426 13268 19432 13320
rect 19484 13268 19490 13320
rect 20622 13268 20628 13320
rect 20680 13308 20686 13320
rect 20958 13311 21016 13317
rect 20958 13308 20970 13311
rect 20680 13280 20970 13308
rect 20680 13268 20686 13280
rect 20958 13277 20970 13280
rect 21004 13308 21016 13311
rect 23492 13308 23520 13407
rect 21004 13280 23520 13308
rect 21004 13277 21016 13280
rect 20958 13271 21016 13277
rect 23658 13268 23664 13320
rect 23716 13268 23722 13320
rect 13357 13243 13415 13249
rect 13357 13209 13369 13243
rect 13403 13240 13415 13243
rect 14139 13243 14197 13249
rect 14139 13240 14151 13243
rect 13403 13212 14151 13240
rect 13403 13209 13415 13212
rect 13357 13203 13415 13209
rect 14139 13209 14151 13212
rect 14185 13209 14197 13243
rect 14139 13203 14197 13209
rect 14737 13243 14795 13249
rect 14737 13209 14749 13243
rect 14783 13240 14795 13243
rect 15289 13243 15347 13249
rect 15289 13240 15301 13243
rect 14783 13212 15301 13240
rect 14783 13209 14795 13212
rect 14737 13203 14795 13209
rect 15289 13209 15301 13212
rect 15335 13209 15347 13243
rect 15289 13203 15347 13209
rect 1578 13132 1584 13184
rect 1636 13132 1642 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7055 13175 7113 13181
rect 7055 13172 7067 13175
rect 6972 13144 7067 13172
rect 6972 13132 6978 13144
rect 7055 13141 7067 13144
rect 7101 13141 7113 13175
rect 7055 13135 7113 13141
rect 15657 13175 15715 13181
rect 15657 13141 15669 13175
rect 15703 13172 15715 13175
rect 15838 13172 15844 13184
rect 15703 13144 15844 13172
rect 15703 13141 15715 13144
rect 15657 13135 15715 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 19208 13144 19257 13172
rect 19208 13132 19214 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 20855 13175 20913 13181
rect 20855 13172 20867 13175
rect 20772 13144 20867 13172
rect 20772 13132 20778 13144
rect 20855 13141 20867 13144
rect 20901 13141 20913 13175
rect 20855 13135 20913 13141
rect 1104 13082 24012 13104
rect 1104 13030 4473 13082
rect 4525 13030 4537 13082
rect 4589 13030 4601 13082
rect 4653 13030 4665 13082
rect 4717 13030 4729 13082
rect 4781 13030 10200 13082
rect 10252 13030 10264 13082
rect 10316 13030 10328 13082
rect 10380 13030 10392 13082
rect 10444 13030 10456 13082
rect 10508 13030 15927 13082
rect 15979 13030 15991 13082
rect 16043 13030 16055 13082
rect 16107 13030 16119 13082
rect 16171 13030 16183 13082
rect 16235 13030 21654 13082
rect 21706 13030 21718 13082
rect 21770 13030 21782 13082
rect 21834 13030 21846 13082
rect 21898 13030 21910 13082
rect 21962 13030 24012 13082
rect 1104 13008 24012 13030
rect 2746 12940 6776 12968
rect 1578 12860 1584 12912
rect 1636 12900 1642 12912
rect 2746 12900 2774 12940
rect 6748 12900 6776 12940
rect 6914 12928 6920 12980
rect 6972 12928 6978 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10229 12971 10287 12977
rect 10229 12968 10241 12971
rect 10008 12940 10241 12968
rect 10008 12928 10014 12940
rect 10229 12937 10241 12940
rect 10275 12937 10287 12971
rect 10229 12931 10287 12937
rect 14090 12928 14096 12980
rect 14148 12968 14154 12980
rect 14369 12971 14427 12977
rect 14369 12968 14381 12971
rect 14148 12940 14381 12968
rect 14148 12928 14154 12940
rect 14369 12937 14381 12940
rect 14415 12937 14427 12971
rect 14369 12931 14427 12937
rect 19150 12928 19156 12980
rect 19208 12928 19214 12980
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12937 20315 12971
rect 20257 12931 20315 12937
rect 8481 12903 8539 12909
rect 8481 12900 8493 12903
rect 1636 12872 2774 12900
rect 5000 12872 5672 12900
rect 6748 12872 8493 12900
rect 1636 12860 1642 12872
rect 5000 12844 5028 12872
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 4408 12835 4466 12841
rect 4408 12801 4420 12835
rect 4454 12832 4466 12835
rect 4798 12832 4804 12844
rect 4454 12804 4804 12832
rect 4454 12801 4466 12804
rect 4408 12795 4466 12801
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 4982 12792 4988 12844
rect 5040 12792 5046 12844
rect 5644 12841 5672 12872
rect 8481 12869 8493 12872
rect 8527 12900 8539 12903
rect 8527 12872 9168 12900
rect 8527 12869 8539 12872
rect 8481 12863 8539 12869
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12832 5135 12835
rect 5491 12835 5549 12841
rect 5491 12832 5503 12835
rect 5123 12804 5503 12832
rect 5123 12801 5135 12804
rect 5077 12795 5135 12801
rect 5491 12801 5503 12804
rect 5537 12801 5549 12835
rect 5491 12795 5549 12801
rect 5594 12835 5672 12841
rect 5594 12801 5606 12835
rect 5640 12804 5672 12835
rect 5640 12801 5652 12804
rect 5594 12795 5652 12801
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 9140 12841 9168 12872
rect 19426 12860 19432 12912
rect 19484 12900 19490 12912
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 19484 12872 19809 12900
rect 19484 12860 19490 12872
rect 19797 12869 19809 12872
rect 19843 12869 19855 12903
rect 19797 12863 19855 12869
rect 19978 12860 19984 12912
rect 20036 12900 20042 12912
rect 20272 12900 20300 12931
rect 20622 12928 20628 12980
rect 20680 12928 20686 12980
rect 20714 12928 20720 12980
rect 20772 12928 20778 12980
rect 20036 12872 20300 12900
rect 20036 12860 20042 12872
rect 8573 12835 8631 12841
rect 8573 12801 8585 12835
rect 8619 12832 8631 12835
rect 8987 12835 9045 12841
rect 8987 12832 8999 12835
rect 8619 12804 8999 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 8987 12801 8999 12804
rect 9033 12801 9045 12835
rect 8987 12795 9045 12801
rect 9090 12835 9168 12841
rect 9090 12801 9102 12835
rect 9136 12804 9168 12835
rect 9136 12801 9148 12804
rect 9090 12795 9148 12801
rect 10410 12792 10416 12844
rect 10468 12792 10474 12844
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12832 10655 12835
rect 10870 12832 10876 12844
rect 10643 12804 10876 12832
rect 10643 12801 10655 12804
rect 10597 12795 10655 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12832 14059 12835
rect 14610 12835 14668 12841
rect 14610 12832 14622 12835
rect 14047 12804 14622 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 14610 12801 14622 12804
rect 14656 12832 14668 12835
rect 14918 12832 14924 12844
rect 14656 12804 14924 12832
rect 14656 12801 14668 12804
rect 14610 12795 14668 12801
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 19245 12835 19303 12841
rect 19245 12801 19257 12835
rect 19291 12832 19303 12835
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19291 12804 19625 12832
rect 19291 12801 19303 12804
rect 19245 12795 19303 12801
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 21234 12835 21292 12841
rect 21234 12801 21246 12835
rect 21280 12832 21292 12835
rect 21358 12832 21364 12844
rect 21280 12804 21364 12832
rect 21280 12801 21292 12804
rect 21234 12795 21292 12801
rect 21358 12792 21364 12804
rect 21416 12832 21422 12844
rect 21416 12804 22094 12832
rect 21416 12792 21422 12804
rect 2746 12736 5120 12764
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 2746 12696 2774 12736
rect 1627 12668 2774 12696
rect 4479 12699 4537 12705
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 4479 12665 4491 12699
rect 4525 12696 4537 12699
rect 4706 12696 4712 12708
rect 4525 12668 4712 12696
rect 4525 12665 4537 12668
rect 4479 12659 4537 12665
rect 4706 12656 4712 12668
rect 4764 12656 4770 12708
rect 5092 12696 5120 12736
rect 5258 12724 5264 12776
rect 5316 12724 5322 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 6914 12764 6920 12776
rect 6871 12736 6920 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 7024 12696 7052 12792
rect 7098 12724 7104 12776
rect 7156 12764 7162 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7156 12736 7849 12764
rect 7156 12724 7162 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 5092 12668 7052 12696
rect 7374 12656 7380 12708
rect 7432 12696 7438 12708
rect 7653 12699 7711 12705
rect 7653 12696 7665 12699
rect 7432 12668 7665 12696
rect 7432 12656 7438 12668
rect 7653 12665 7665 12668
rect 7699 12665 7711 12699
rect 7653 12659 7711 12665
rect 4338 12588 4344 12640
rect 4396 12628 4402 12640
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 4396 12600 4629 12628
rect 4396 12588 4402 12600
rect 4617 12597 4629 12600
rect 4663 12597 4675 12631
rect 7852 12628 7880 12727
rect 8662 12724 8668 12776
rect 8720 12724 8726 12776
rect 13814 12724 13820 12776
rect 13872 12724 13878 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12764 13967 12767
rect 14507 12767 14565 12773
rect 14507 12764 14519 12767
rect 13955 12736 14519 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 14507 12733 14519 12736
rect 14553 12733 14565 12767
rect 14507 12727 14565 12733
rect 19058 12724 19064 12776
rect 19116 12764 19122 12776
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 19116 12736 19349 12764
rect 19116 12724 19122 12736
rect 19337 12733 19349 12736
rect 19383 12733 19395 12767
rect 19337 12727 19395 12733
rect 20809 12767 20867 12773
rect 20809 12733 20821 12767
rect 20855 12733 20867 12767
rect 22066 12764 22094 12804
rect 23382 12792 23388 12844
rect 23440 12832 23446 12844
rect 23661 12835 23719 12841
rect 23661 12832 23673 12835
rect 23440 12804 23673 12832
rect 23440 12792 23446 12804
rect 23661 12801 23673 12804
rect 23707 12801 23719 12835
rect 23661 12795 23719 12801
rect 22066 12736 23520 12764
rect 20809 12727 20867 12733
rect 8021 12699 8079 12705
rect 8021 12665 8033 12699
rect 8067 12696 8079 12699
rect 8294 12696 8300 12708
rect 8067 12668 8300 12696
rect 8067 12665 8079 12668
rect 8021 12659 8079 12665
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 17034 12656 17040 12708
rect 17092 12696 17098 12708
rect 20824 12696 20852 12727
rect 23198 12696 23204 12708
rect 17092 12668 23204 12696
rect 17092 12656 17098 12668
rect 23198 12656 23204 12668
rect 23256 12656 23262 12708
rect 23492 12705 23520 12736
rect 23477 12699 23535 12705
rect 23477 12665 23489 12699
rect 23523 12665 23535 12699
rect 23477 12659 23535 12665
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 7852 12600 8125 12628
rect 4617 12591 4675 12597
rect 8113 12597 8125 12600
rect 8159 12597 8171 12631
rect 8113 12591 8171 12597
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 11054 12628 11060 12640
rect 8260 12600 11060 12628
rect 8260 12588 8266 12600
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 18230 12588 18236 12640
rect 18288 12628 18294 12640
rect 18785 12631 18843 12637
rect 18785 12628 18797 12631
rect 18288 12600 18797 12628
rect 18288 12588 18294 12600
rect 18785 12597 18797 12600
rect 18831 12597 18843 12631
rect 18785 12591 18843 12597
rect 20898 12588 20904 12640
rect 20956 12628 20962 12640
rect 21131 12631 21189 12637
rect 21131 12628 21143 12631
rect 20956 12600 21143 12628
rect 20956 12588 20962 12600
rect 21131 12597 21143 12600
rect 21177 12597 21189 12631
rect 21131 12591 21189 12597
rect 1104 12538 24012 12560
rect 1104 12486 3813 12538
rect 3865 12486 3877 12538
rect 3929 12486 3941 12538
rect 3993 12486 4005 12538
rect 4057 12486 4069 12538
rect 4121 12486 9540 12538
rect 9592 12486 9604 12538
rect 9656 12486 9668 12538
rect 9720 12486 9732 12538
rect 9784 12486 9796 12538
rect 9848 12486 15267 12538
rect 15319 12486 15331 12538
rect 15383 12486 15395 12538
rect 15447 12486 15459 12538
rect 15511 12486 15523 12538
rect 15575 12486 20994 12538
rect 21046 12486 21058 12538
rect 21110 12486 21122 12538
rect 21174 12486 21186 12538
rect 21238 12486 21250 12538
rect 21302 12486 24012 12538
rect 1104 12464 24012 12486
rect 5350 12424 5356 12436
rect 4632 12396 5356 12424
rect 4632 12297 4660 12396
rect 5350 12384 5356 12396
rect 5408 12424 5414 12436
rect 6914 12424 6920 12436
rect 5408 12396 6920 12424
rect 5408 12384 5414 12396
rect 6914 12384 6920 12396
rect 6972 12424 6978 12436
rect 7282 12424 7288 12436
rect 6972 12396 7288 12424
rect 6972 12384 6978 12396
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 10410 12424 10416 12436
rect 9723 12396 10416 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 6825 12359 6883 12365
rect 6825 12325 6837 12359
rect 6871 12356 6883 12359
rect 7374 12356 7380 12368
rect 6871 12328 7380 12356
rect 6871 12325 6883 12328
rect 6825 12319 6883 12325
rect 4617 12291 4675 12297
rect 4617 12257 4629 12291
rect 4663 12257 4675 12291
rect 4617 12251 4675 12257
rect 4706 12248 4712 12300
rect 4764 12248 4770 12300
rect 6932 12229 6960 12328
rect 7374 12316 7380 12328
rect 7432 12316 7438 12368
rect 10781 12359 10839 12365
rect 10781 12356 10793 12359
rect 9508 12328 10793 12356
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12288 8079 12291
rect 8202 12288 8208 12300
rect 8067 12260 8208 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12288 8723 12291
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 8711 12260 9321 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9309 12251 9367 12257
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12189 6699 12223
rect 6641 12183 6699 12189
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 6656 12152 6684 12183
rect 7098 12180 7104 12232
rect 7156 12180 7162 12232
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12220 7343 12223
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7331 12192 7849 12220
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8294 12180 8300 12232
rect 8352 12180 8358 12232
rect 7116 12152 7144 12180
rect 7745 12155 7803 12161
rect 7745 12152 7757 12155
rect 6656 12124 7144 12152
rect 7208 12124 7757 12152
rect 4798 12044 4804 12096
rect 4856 12044 4862 12096
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5534 12084 5540 12096
rect 5215 12056 5540 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 6457 12087 6515 12093
rect 6457 12053 6469 12087
rect 6503 12084 6515 12087
rect 7208 12084 7236 12124
rect 7745 12121 7757 12124
rect 7791 12121 7803 12155
rect 7745 12115 7803 12121
rect 8478 12112 8484 12164
rect 8536 12112 8542 12164
rect 9324 12152 9352 12251
rect 9508 12229 9536 12328
rect 10060 12297 10088 12328
rect 10781 12325 10793 12328
rect 10827 12325 10839 12359
rect 19889 12359 19947 12365
rect 10781 12319 10839 12325
rect 11164 12328 11836 12356
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12257 10379 12291
rect 10321 12251 10379 12257
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 9968 12152 9996 12183
rect 9324 12124 9996 12152
rect 10042 12112 10048 12164
rect 10100 12152 10106 12164
rect 10336 12152 10364 12251
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12220 10471 12223
rect 10594 12220 10600 12232
rect 10459 12192 10600 12220
rect 10459 12189 10471 12192
rect 10413 12183 10471 12189
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 11164 12229 11192 12328
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12257 11299 12291
rect 11241 12251 11299 12257
rect 11149 12223 11207 12229
rect 11149 12189 11161 12223
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 10100 12124 10364 12152
rect 11256 12152 11284 12251
rect 11606 12152 11612 12164
rect 11256 12124 11612 12152
rect 10100 12112 10106 12124
rect 11606 12112 11612 12124
rect 11664 12112 11670 12164
rect 11808 12161 11836 12328
rect 19889 12325 19901 12359
rect 19935 12356 19947 12359
rect 19978 12356 19984 12368
rect 19935 12328 19984 12356
rect 19935 12325 19947 12328
rect 19889 12319 19947 12325
rect 15562 12248 15568 12300
rect 15620 12288 15626 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15620 12260 15669 12288
rect 15620 12248 15626 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 16025 12291 16083 12297
rect 16025 12257 16037 12291
rect 16071 12288 16083 12291
rect 16482 12288 16488 12300
rect 16071 12260 16488 12288
rect 16071 12257 16083 12260
rect 16025 12251 16083 12257
rect 16482 12248 16488 12260
rect 16540 12248 16546 12300
rect 18966 12248 18972 12300
rect 19024 12288 19030 12300
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 19024 12260 19257 12288
rect 19024 12248 19030 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19521 12291 19579 12297
rect 19521 12288 19533 12291
rect 19484 12260 19533 12288
rect 19484 12248 19490 12260
rect 19521 12257 19533 12260
rect 19567 12257 19579 12291
rect 19521 12251 19579 12257
rect 12494 12223 12552 12229
rect 12494 12189 12506 12223
rect 12540 12220 12552 12223
rect 12618 12220 12624 12232
rect 12540 12192 12624 12220
rect 12540 12189 12552 12192
rect 12494 12183 12552 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15804 12192 15853 12220
rect 15804 12180 15810 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 16368 12223 16426 12229
rect 16368 12189 16380 12223
rect 16414 12220 16426 12223
rect 17034 12220 17040 12232
rect 16414 12192 17040 12220
rect 16414 12189 16426 12192
rect 16368 12183 16426 12189
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 11793 12155 11851 12161
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 11882 12152 11888 12164
rect 11839 12124 11888 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 19536 12152 19564 12251
rect 19613 12223 19671 12229
rect 19613 12189 19625 12223
rect 19659 12220 19671 12223
rect 19904 12220 19932 12319
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 20898 12248 20904 12300
rect 20956 12248 20962 12300
rect 21085 12291 21143 12297
rect 21085 12257 21097 12291
rect 21131 12288 21143 12291
rect 22186 12288 22192 12300
rect 21131 12260 22192 12288
rect 21131 12257 21143 12260
rect 21085 12251 21143 12257
rect 22186 12248 22192 12260
rect 22244 12248 22250 12300
rect 19659 12192 19932 12220
rect 20073 12223 20131 12229
rect 19659 12189 19671 12192
rect 19613 12183 19671 12189
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12220 20867 12223
rect 21358 12220 21364 12232
rect 20855 12192 21364 12220
rect 20855 12189 20867 12192
rect 20809 12183 20867 12189
rect 20088 12152 20116 12183
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 19536 12124 20484 12152
rect 6503 12056 7236 12084
rect 6503 12053 6515 12056
rect 6457 12047 6515 12053
rect 7374 12044 7380 12096
rect 7432 12044 7438 12096
rect 11422 12044 11428 12096
rect 11480 12044 11486 12096
rect 12434 12093 12440 12096
rect 12391 12087 12440 12093
rect 12391 12053 12403 12087
rect 12437 12053 12440 12087
rect 12391 12047 12440 12053
rect 12434 12044 12440 12047
rect 12492 12044 12498 12096
rect 16439 12087 16497 12093
rect 16439 12053 16451 12087
rect 16485 12084 16497 12087
rect 17126 12084 17132 12096
rect 16485 12056 17132 12084
rect 16485 12053 16497 12056
rect 16439 12047 16497 12053
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 20456 12093 20484 12124
rect 20257 12087 20315 12093
rect 20257 12084 20269 12087
rect 20220 12056 20269 12084
rect 20220 12044 20226 12056
rect 20257 12053 20269 12056
rect 20303 12053 20315 12087
rect 20257 12047 20315 12053
rect 20441 12087 20499 12093
rect 20441 12053 20453 12087
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 1104 11994 24012 12016
rect 1104 11942 4473 11994
rect 4525 11942 4537 11994
rect 4589 11942 4601 11994
rect 4653 11942 4665 11994
rect 4717 11942 4729 11994
rect 4781 11942 10200 11994
rect 10252 11942 10264 11994
rect 10316 11942 10328 11994
rect 10380 11942 10392 11994
rect 10444 11942 10456 11994
rect 10508 11942 15927 11994
rect 15979 11942 15991 11994
rect 16043 11942 16055 11994
rect 16107 11942 16119 11994
rect 16171 11942 16183 11994
rect 16235 11942 21654 11994
rect 21706 11942 21718 11994
rect 21770 11942 21782 11994
rect 21834 11942 21846 11994
rect 21898 11942 21910 11994
rect 21962 11942 24012 11994
rect 1104 11920 24012 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 4798 11880 4804 11892
rect 1627 11852 4804 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 8478 11880 8484 11892
rect 8343 11852 8484 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 10100 11852 10241 11880
rect 10100 11840 10106 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 10229 11843 10287 11849
rect 10321 11883 10379 11889
rect 10321 11849 10333 11883
rect 10367 11880 10379 11883
rect 10594 11880 10600 11892
rect 10367 11852 10600 11880
rect 10367 11849 10379 11852
rect 10321 11843 10379 11849
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 10870 11840 10876 11892
rect 10928 11840 10934 11892
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 13814 11880 13820 11892
rect 12860 11852 13820 11880
rect 12860 11840 12866 11852
rect 13814 11840 13820 11852
rect 13872 11880 13878 11892
rect 13872 11852 16804 11880
rect 13872 11840 13878 11852
rect 3789 11815 3847 11821
rect 3789 11781 3801 11815
rect 3835 11812 3847 11815
rect 5077 11815 5135 11821
rect 5077 11812 5089 11815
rect 3835 11784 5089 11812
rect 3835 11781 3847 11784
rect 3789 11775 3847 11781
rect 5077 11781 5089 11784
rect 5123 11781 5135 11815
rect 5077 11775 5135 11781
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 8202 11812 8208 11824
rect 5500 11784 8208 11812
rect 5500 11772 5506 11784
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 12529 11815 12587 11821
rect 12529 11781 12541 11815
rect 12575 11812 12587 11815
rect 12575 11784 13216 11812
rect 12575 11781 12587 11784
rect 12529 11775 12587 11781
rect 842 11704 848 11756
rect 900 11744 906 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 900 11716 1409 11744
rect 900 11704 906 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 4154 11744 4160 11756
rect 4019 11716 4160 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4264 11608 4292 11707
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4396 11716 4445 11744
rect 4396 11704 4402 11716
rect 4433 11713 4445 11716
rect 4479 11744 4491 11747
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 4479 11716 5733 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 5721 11713 5733 11716
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 7466 11704 7472 11756
rect 7524 11704 7530 11756
rect 13188 11753 13216 11784
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 13035 11747 13093 11753
rect 13035 11744 13047 11747
rect 12667 11716 13047 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 13035 11713 13047 11716
rect 13081 11713 13093 11747
rect 13035 11707 13093 11713
rect 13138 11747 13216 11753
rect 13138 11713 13150 11747
rect 13184 11713 13216 11747
rect 13138 11707 13216 11713
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11676 4675 11679
rect 5169 11679 5227 11685
rect 5169 11676 5181 11679
rect 4663 11648 5181 11676
rect 4663 11645 4675 11648
rect 4617 11639 4675 11645
rect 5169 11645 5181 11648
rect 5215 11645 5227 11679
rect 5169 11639 5227 11645
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 5442 11676 5448 11688
rect 5399 11648 5448 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5534 11636 5540 11688
rect 5592 11636 5598 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7377 11679 7435 11685
rect 7377 11676 7389 11679
rect 7156 11648 7389 11676
rect 7156 11636 7162 11648
rect 7377 11645 7389 11648
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11645 8171 11679
rect 8113 11639 8171 11645
rect 5552 11608 5580 11636
rect 4203 11580 5580 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4632 11552 4660 11580
rect 7742 11568 7748 11620
rect 7800 11608 7806 11620
rect 7929 11611 7987 11617
rect 7929 11608 7941 11611
rect 7800 11580 7941 11608
rect 7800 11568 7806 11580
rect 7929 11577 7941 11580
rect 7975 11577 7987 11611
rect 7929 11571 7987 11577
rect 4614 11500 4620 11552
rect 4672 11500 4678 11552
rect 4709 11543 4767 11549
rect 4709 11509 4721 11543
rect 4755 11540 4767 11543
rect 4982 11540 4988 11552
rect 4755 11512 4988 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5810 11500 5816 11552
rect 5868 11540 5874 11552
rect 5905 11543 5963 11549
rect 5905 11540 5917 11543
rect 5868 11512 5917 11540
rect 5868 11500 5874 11512
rect 5905 11509 5917 11512
rect 5951 11509 5963 11543
rect 5905 11503 5963 11509
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 7837 11543 7895 11549
rect 7837 11540 7849 11543
rect 7708 11512 7849 11540
rect 7708 11500 7714 11512
rect 7837 11509 7849 11512
rect 7883 11540 7895 11543
rect 8128 11540 8156 11639
rect 10502 11636 10508 11688
rect 10560 11636 10566 11688
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11606 11676 11612 11688
rect 11103 11648 11612 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 11606 11636 11612 11648
rect 11664 11676 11670 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11664 11648 11713 11676
rect 11664 11636 11670 11648
rect 11701 11645 11713 11648
rect 11747 11676 11759 11679
rect 11747 11648 12204 11676
rect 11747 11645 11759 11648
rect 11701 11639 11759 11645
rect 11241 11611 11299 11617
rect 11241 11577 11253 11611
rect 11287 11608 11299 11611
rect 11882 11608 11888 11620
rect 11287 11580 11888 11608
rect 11287 11577 11299 11580
rect 11241 11571 11299 11577
rect 11882 11568 11888 11580
rect 11940 11568 11946 11620
rect 12176 11617 12204 11648
rect 12802 11636 12808 11688
rect 12860 11636 12866 11688
rect 13188 11676 13216 11707
rect 15562 11704 15568 11756
rect 15620 11704 15626 11756
rect 15746 11744 15752 11756
rect 15672 11716 15752 11744
rect 15672 11685 15700 11716
rect 15746 11704 15752 11716
rect 15804 11744 15810 11756
rect 15804 11716 16712 11744
rect 15804 11704 15810 11716
rect 13096 11648 13216 11676
rect 15657 11679 15715 11685
rect 13096 11620 13124 11648
rect 15657 11645 15669 11679
rect 15703 11645 15715 11679
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 15657 11639 15715 11645
rect 15948 11648 16221 11676
rect 12161 11611 12219 11617
rect 12161 11577 12173 11611
rect 12207 11577 12219 11611
rect 12161 11571 12219 11577
rect 13078 11568 13084 11620
rect 13136 11568 13142 11620
rect 15948 11552 15976 11648
rect 16209 11645 16221 11648
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 16022 11568 16028 11620
rect 16080 11568 16086 11620
rect 16684 11617 16712 11716
rect 16776 11676 16804 11852
rect 17126 11840 17132 11892
rect 17184 11840 17190 11892
rect 23477 11883 23535 11889
rect 23477 11880 23489 11883
rect 18524 11852 23489 11880
rect 17034 11772 17040 11824
rect 17092 11812 17098 11824
rect 18524 11812 18552 11852
rect 23477 11849 23489 11852
rect 23523 11849 23535 11883
rect 23477 11843 23535 11849
rect 17092 11784 18552 11812
rect 17092 11772 17098 11784
rect 20162 11772 20168 11824
rect 20220 11772 20226 11824
rect 18506 11704 18512 11756
rect 18564 11704 18570 11756
rect 18966 11744 18972 11756
rect 18616 11716 18972 11744
rect 18616 11685 18644 11716
rect 18966 11704 18972 11716
rect 19024 11704 19030 11756
rect 19153 11747 19211 11753
rect 19153 11713 19165 11747
rect 19199 11744 19211 11747
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19199 11716 19993 11744
rect 19199 11713 19211 11716
rect 19153 11707 19211 11713
rect 19981 11713 19993 11716
rect 20027 11713 20039 11747
rect 19981 11707 20039 11713
rect 23658 11704 23664 11756
rect 23716 11704 23722 11756
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 16776 11648 17233 11676
rect 17221 11645 17233 11648
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 18601 11679 18659 11685
rect 18601 11645 18613 11679
rect 18647 11645 18659 11679
rect 18601 11639 18659 11645
rect 16669 11611 16727 11617
rect 16669 11577 16681 11611
rect 16715 11577 16727 11611
rect 16669 11571 16727 11577
rect 18506 11568 18512 11620
rect 18564 11608 18570 11620
rect 18785 11611 18843 11617
rect 18785 11608 18797 11611
rect 18564 11580 18797 11608
rect 18564 11568 18570 11580
rect 18785 11577 18797 11580
rect 18831 11577 18843 11611
rect 18785 11571 18843 11577
rect 7883 11512 8156 11540
rect 9861 11543 9919 11549
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10042 11540 10048 11552
rect 9907 11512 10048 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 11514 11500 11520 11552
rect 11572 11500 11578 11552
rect 15930 11500 15936 11552
rect 15988 11500 15994 11552
rect 16390 11500 16396 11552
rect 16448 11500 16454 11552
rect 18141 11543 18199 11549
rect 18141 11509 18153 11543
rect 18187 11540 18199 11543
rect 18414 11540 18420 11552
rect 18187 11512 18420 11540
rect 18187 11509 18199 11512
rect 18141 11503 18199 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 19797 11543 19855 11549
rect 19797 11509 19809 11543
rect 19843 11540 19855 11543
rect 20714 11540 20720 11552
rect 19843 11512 20720 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 1104 11450 24012 11472
rect 1104 11398 3813 11450
rect 3865 11398 3877 11450
rect 3929 11398 3941 11450
rect 3993 11398 4005 11450
rect 4057 11398 4069 11450
rect 4121 11398 9540 11450
rect 9592 11398 9604 11450
rect 9656 11398 9668 11450
rect 9720 11398 9732 11450
rect 9784 11398 9796 11450
rect 9848 11398 15267 11450
rect 15319 11398 15331 11450
rect 15383 11398 15395 11450
rect 15447 11398 15459 11450
rect 15511 11398 15523 11450
rect 15575 11398 20994 11450
rect 21046 11398 21058 11450
rect 21110 11398 21122 11450
rect 21174 11398 21186 11450
rect 21238 11398 21250 11450
rect 21302 11398 24012 11450
rect 1104 11376 24012 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 4890 11336 4896 11348
rect 1627 11308 4896 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 11054 11336 11060 11348
rect 10560 11308 11060 11336
rect 10560 11296 10566 11308
rect 11054 11296 11060 11308
rect 11112 11336 11118 11348
rect 11112 11308 11744 11336
rect 11112 11296 11118 11308
rect 9306 11228 9312 11280
rect 9364 11268 9370 11280
rect 9585 11271 9643 11277
rect 9585 11268 9597 11271
rect 9364 11240 9597 11268
rect 9364 11228 9370 11240
rect 9585 11237 9597 11240
rect 9631 11237 9643 11271
rect 11149 11271 11207 11277
rect 11149 11268 11161 11271
rect 9585 11231 9643 11237
rect 9968 11240 11161 11268
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4801 11203 4859 11209
rect 4801 11200 4813 11203
rect 4396 11172 4813 11200
rect 4396 11160 4402 11172
rect 4801 11169 4813 11172
rect 4847 11169 4859 11203
rect 4801 11163 4859 11169
rect 5074 11160 5080 11212
rect 5132 11160 5138 11212
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 5491 11172 6914 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 4614 11092 4620 11144
rect 4672 11132 4678 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 4672 11104 4721 11132
rect 4672 11092 4678 11104
rect 4709 11101 4721 11104
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 5810 11092 5816 11144
rect 5868 11092 5874 11144
rect 6886 11132 6914 11172
rect 7650 11160 7656 11212
rect 7708 11160 7714 11212
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 7929 11203 7987 11209
rect 7929 11200 7941 11203
rect 7892 11172 7941 11200
rect 7892 11160 7898 11172
rect 7929 11169 7941 11172
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 6886 11104 7573 11132
rect 7561 11101 7573 11104
rect 7607 11132 7619 11135
rect 7742 11132 7748 11144
rect 7607 11104 7748 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 9968 11141 9996 11240
rect 11149 11237 11161 11240
rect 11195 11237 11207 11271
rect 11149 11231 11207 11237
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 5626 11024 5632 11076
rect 5684 11024 5690 11076
rect 8570 11024 8576 11076
rect 8628 11064 8634 11076
rect 10152 11064 10180 11163
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 11716 11209 11744 11308
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 11940 11308 11989 11336
rect 11940 11296 11946 11308
rect 11977 11305 11989 11308
rect 12023 11305 12035 11339
rect 11977 11299 12035 11305
rect 14921 11339 14979 11345
rect 14921 11305 14933 11339
rect 14967 11336 14979 11339
rect 15286 11336 15292 11348
rect 14967 11308 15292 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15286 11296 15292 11308
rect 15344 11336 15350 11348
rect 15654 11336 15660 11348
rect 15344 11308 15660 11336
rect 15344 11296 15350 11308
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16853 11339 16911 11345
rect 16853 11305 16865 11339
rect 16899 11336 16911 11339
rect 18506 11336 18512 11348
rect 16899 11308 18512 11336
rect 16899 11305 16911 11308
rect 16853 11299 16911 11305
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 23477 11271 23535 11277
rect 23477 11268 23489 11271
rect 12400 11240 12664 11268
rect 12400 11228 12406 11240
rect 11609 11203 11667 11209
rect 11609 11200 11621 11203
rect 11480 11172 11621 11200
rect 11480 11160 11486 11172
rect 11609 11169 11621 11172
rect 11655 11169 11667 11203
rect 11609 11163 11667 11169
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 12434 11160 12440 11212
rect 12492 11160 12498 11212
rect 12636 11209 12664 11240
rect 15764 11240 23489 11268
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11200 12679 11203
rect 13262 11200 13268 11212
rect 12667 11172 13268 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 13262 11160 13268 11172
rect 13320 11200 13326 11212
rect 14277 11203 14335 11209
rect 14277 11200 14289 11203
rect 13320 11172 14289 11200
rect 13320 11160 13326 11172
rect 14277 11169 14289 11172
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 11514 11092 11520 11144
rect 11572 11092 11578 11144
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 15151 11135 15209 11141
rect 15151 11132 15163 11135
rect 14599 11104 15163 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 15151 11101 15163 11104
rect 15197 11132 15209 11135
rect 15764 11132 15792 11240
rect 23477 11237 23489 11240
rect 23523 11237 23535 11271
rect 23477 11231 23535 11237
rect 15930 11160 15936 11212
rect 15988 11160 15994 11212
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 16298 11200 16304 11212
rect 16255 11172 16304 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 18380 11172 18429 11200
rect 18380 11160 18386 11172
rect 18417 11169 18429 11172
rect 18463 11200 18475 11203
rect 19242 11200 19248 11212
rect 18463 11172 19248 11200
rect 18463 11169 18475 11172
rect 18417 11163 18475 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11200 22155 11203
rect 22646 11200 22652 11212
rect 22143 11172 22652 11200
rect 22143 11169 22155 11172
rect 22097 11163 22155 11169
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 15197 11104 15792 11132
rect 15197 11101 15209 11104
rect 15151 11095 15209 11101
rect 15838 11092 15844 11144
rect 15896 11092 15902 11144
rect 16390 11092 16396 11144
rect 16448 11132 16454 11144
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 16448 11104 16681 11132
rect 16448 11092 16454 11104
rect 16669 11101 16681 11104
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 18230 11092 18236 11144
rect 18288 11092 18294 11144
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 21913 11135 21971 11141
rect 21913 11132 21925 11135
rect 21600 11104 21925 11132
rect 21600 11092 21606 11104
rect 21913 11101 21925 11104
rect 21959 11101 21971 11135
rect 21913 11095 21971 11101
rect 22982 11135 23040 11141
rect 22982 11101 22994 11135
rect 23028 11132 23040 11135
rect 23290 11132 23296 11144
rect 23028 11104 23296 11132
rect 23028 11101 23040 11104
rect 22982 11095 23040 11101
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 23382 11092 23388 11144
rect 23440 11132 23446 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 23440 11104 23673 11132
rect 23440 11092 23446 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 8628 11036 10180 11064
rect 12345 11067 12403 11073
rect 8628 11024 8634 11036
rect 12345 11033 12357 11067
rect 12391 11064 12403 11067
rect 12618 11064 12624 11076
rect 12391 11036 12624 11064
rect 12391 11033 12403 11036
rect 12345 11027 12403 11033
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 14461 11067 14519 11073
rect 14461 11033 14473 11067
rect 14507 11064 14519 11067
rect 15059 11067 15117 11073
rect 15059 11064 15071 11067
rect 14507 11036 15071 11064
rect 14507 11033 14519 11036
rect 14461 11027 14519 11033
rect 15059 11033 15071 11036
rect 15105 11033 15117 11067
rect 15059 11027 15117 11033
rect 16482 11024 16488 11076
rect 16540 11024 16546 11076
rect 21269 11067 21327 11073
rect 21269 11033 21281 11067
rect 21315 11064 21327 11067
rect 21358 11064 21364 11076
rect 21315 11036 21364 11064
rect 21315 11033 21327 11036
rect 21269 11027 21327 11033
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 21450 11024 21456 11076
rect 21508 11024 21514 11076
rect 21637 11067 21695 11073
rect 21637 11033 21649 11067
rect 21683 11064 21695 11067
rect 21729 11067 21787 11073
rect 21729 11064 21741 11067
rect 21683 11036 21741 11064
rect 21683 11033 21695 11036
rect 21637 11027 21695 11033
rect 21729 11033 21741 11036
rect 21775 11033 21787 11067
rect 21729 11027 21787 11033
rect 17678 10956 17684 11008
rect 17736 10996 17742 11008
rect 17865 10999 17923 11005
rect 17865 10996 17877 10999
rect 17736 10968 17877 10996
rect 17736 10956 17742 10968
rect 17865 10965 17877 10968
rect 17911 10965 17923 10999
rect 17865 10959 17923 10965
rect 18322 10956 18328 11008
rect 18380 10956 18386 11008
rect 22879 10999 22937 11005
rect 22879 10965 22891 10999
rect 22925 10996 22937 10999
rect 23014 10996 23020 11008
rect 22925 10968 23020 10996
rect 22925 10965 22937 10968
rect 22879 10959 22937 10965
rect 23014 10956 23020 10968
rect 23072 10956 23078 11008
rect 1104 10906 24012 10928
rect 1104 10854 4473 10906
rect 4525 10854 4537 10906
rect 4589 10854 4601 10906
rect 4653 10854 4665 10906
rect 4717 10854 4729 10906
rect 4781 10854 10200 10906
rect 10252 10854 10264 10906
rect 10316 10854 10328 10906
rect 10380 10854 10392 10906
rect 10444 10854 10456 10906
rect 10508 10854 15927 10906
rect 15979 10854 15991 10906
rect 16043 10854 16055 10906
rect 16107 10854 16119 10906
rect 16171 10854 16183 10906
rect 16235 10854 21654 10906
rect 21706 10854 21718 10906
rect 21770 10854 21782 10906
rect 21834 10854 21846 10906
rect 21898 10854 21910 10906
rect 21962 10854 24012 10906
rect 1104 10832 24012 10854
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 5813 10795 5871 10801
rect 5813 10792 5825 10795
rect 5684 10764 5825 10792
rect 5684 10752 5690 10764
rect 5813 10761 5825 10764
rect 5859 10761 5871 10795
rect 5813 10755 5871 10761
rect 13357 10795 13415 10801
rect 13357 10761 13369 10795
rect 13403 10792 13415 10795
rect 13722 10792 13728 10804
rect 13403 10764 13728 10792
rect 13403 10761 13415 10764
rect 13357 10755 13415 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10761 13875 10795
rect 13817 10755 13875 10761
rect 14001 10795 14059 10801
rect 14001 10761 14013 10795
rect 14047 10792 14059 10795
rect 18049 10795 18107 10801
rect 14047 10764 14320 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 13538 10684 13544 10736
rect 13596 10684 13602 10736
rect 13832 10724 13860 10755
rect 13832 10696 14228 10724
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 4798 10656 4804 10668
rect 1627 10628 4804 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5000 10520 5028 10619
rect 13170 10616 13176 10668
rect 13228 10616 13234 10668
rect 13262 10616 13268 10668
rect 13320 10616 13326 10668
rect 13556 10656 13584 10684
rect 13633 10659 13691 10665
rect 13633 10656 13645 10659
rect 13556 10628 13645 10656
rect 13633 10625 13645 10628
rect 13679 10625 13691 10659
rect 13633 10619 13691 10625
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5132 10560 5641 10588
rect 5132 10548 5138 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 13538 10548 13544 10600
rect 13596 10548 13602 10600
rect 5442 10520 5448 10532
rect 5000 10492 5448 10520
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 13449 10523 13507 10529
rect 13449 10489 13461 10523
rect 13495 10520 13507 10523
rect 14108 10520 14136 10619
rect 13495 10492 14136 10520
rect 14200 10520 14228 10696
rect 14292 10665 14320 10764
rect 18049 10761 18061 10795
rect 18095 10792 18107 10795
rect 18322 10792 18328 10804
rect 18095 10764 18328 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 18414 10752 18420 10804
rect 18472 10752 18478 10804
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 18690 10792 18696 10804
rect 18555 10764 18696 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 15286 10684 15292 10736
rect 15344 10684 15350 10736
rect 15473 10727 15531 10733
rect 15473 10693 15485 10727
rect 15519 10724 15531 10727
rect 15746 10724 15752 10736
rect 15519 10696 15752 10724
rect 15519 10693 15531 10696
rect 15473 10687 15531 10693
rect 15746 10684 15752 10696
rect 15804 10724 15810 10736
rect 23017 10727 23075 10733
rect 15804 10696 15976 10724
rect 15804 10684 15810 10696
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 15304 10588 15332 10684
rect 15948 10665 15976 10696
rect 19168 10696 22416 10724
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 19168 10600 19196 10696
rect 20714 10616 20720 10668
rect 20772 10616 20778 10668
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10656 21511 10659
rect 21634 10656 21640 10668
rect 21499 10628 21640 10656
rect 21499 10625 21511 10628
rect 21453 10619 21511 10625
rect 21634 10616 21640 10628
rect 21692 10616 21698 10668
rect 22094 10616 22100 10668
rect 22152 10656 22158 10668
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 22152 10628 22201 10656
rect 22152 10616 22158 10628
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 15749 10591 15807 10597
rect 15749 10588 15761 10591
rect 15304 10560 15761 10588
rect 15749 10557 15761 10560
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 18693 10591 18751 10597
rect 18693 10557 18705 10591
rect 18739 10588 18751 10591
rect 19150 10588 19156 10600
rect 18739 10560 19156 10588
rect 18739 10557 18751 10560
rect 18693 10551 18751 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 20898 10588 20904 10600
rect 20855 10560 20904 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 20898 10548 20904 10560
rect 20956 10588 20962 10600
rect 21085 10591 21143 10597
rect 21085 10588 21097 10591
rect 20956 10560 21097 10588
rect 20956 10548 20962 10560
rect 21085 10557 21097 10560
rect 21131 10557 21143 10591
rect 21085 10551 21143 10557
rect 21542 10548 21548 10600
rect 21600 10548 21606 10600
rect 22002 10548 22008 10600
rect 22060 10588 22066 10600
rect 22388 10597 22416 10696
rect 23017 10693 23029 10727
rect 23063 10724 23075 10727
rect 23063 10696 23704 10724
rect 23063 10693 23075 10696
rect 23017 10687 23075 10693
rect 23676 10665 23704 10696
rect 23109 10659 23167 10665
rect 23109 10625 23121 10659
rect 23155 10656 23167 10659
rect 23523 10659 23581 10665
rect 23523 10656 23535 10659
rect 23155 10628 23535 10656
rect 23155 10625 23167 10628
rect 23109 10619 23167 10625
rect 23523 10625 23535 10628
rect 23569 10625 23581 10659
rect 23523 10619 23581 10625
rect 23626 10659 23704 10665
rect 23626 10625 23638 10659
rect 23672 10656 23704 10659
rect 23672 10628 24072 10656
rect 23672 10625 23684 10628
rect 23626 10619 23684 10625
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22060 10560 22293 10588
rect 22060 10548 22066 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 22373 10591 22431 10597
rect 22373 10557 22385 10591
rect 22419 10557 22431 10591
rect 22373 10551 22431 10557
rect 23198 10548 23204 10600
rect 23256 10548 23262 10600
rect 15930 10520 15936 10532
rect 14200 10492 15936 10520
rect 13495 10489 13507 10492
rect 13449 10483 13507 10489
rect 15930 10480 15936 10492
rect 15988 10480 15994 10532
rect 19610 10480 19616 10532
rect 19668 10520 19674 10532
rect 21821 10523 21879 10529
rect 21821 10520 21833 10523
rect 19668 10492 21833 10520
rect 19668 10480 19674 10492
rect 21821 10489 21833 10492
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 842 10412 848 10464
rect 900 10452 906 10464
rect 1397 10455 1455 10461
rect 1397 10452 1409 10455
rect 900 10424 1409 10452
rect 900 10412 906 10424
rect 1397 10421 1409 10424
rect 1443 10421 1455 10455
rect 1397 10415 1455 10421
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 5353 10455 5411 10461
rect 5353 10452 5365 10455
rect 5316 10424 5365 10452
rect 5316 10412 5322 10424
rect 5353 10421 5365 10424
rect 5399 10421 5411 10455
rect 5353 10415 5411 10421
rect 14274 10412 14280 10464
rect 14332 10412 14338 10464
rect 15657 10455 15715 10461
rect 15657 10421 15669 10455
rect 15703 10452 15715 10455
rect 15838 10452 15844 10464
rect 15703 10424 15844 10452
rect 15703 10421 15715 10424
rect 15657 10415 15715 10421
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 16114 10412 16120 10464
rect 16172 10412 16178 10464
rect 19978 10412 19984 10464
rect 20036 10412 20042 10464
rect 20349 10455 20407 10461
rect 20349 10421 20361 10455
rect 20395 10452 20407 10455
rect 20438 10452 20444 10464
rect 20395 10424 20444 10452
rect 20395 10421 20407 10424
rect 20349 10415 20407 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 22646 10412 22652 10464
rect 22704 10412 22710 10464
rect 1104 10362 24012 10384
rect 1104 10310 3813 10362
rect 3865 10310 3877 10362
rect 3929 10310 3941 10362
rect 3993 10310 4005 10362
rect 4057 10310 4069 10362
rect 4121 10310 9540 10362
rect 9592 10310 9604 10362
rect 9656 10310 9668 10362
rect 9720 10310 9732 10362
rect 9784 10310 9796 10362
rect 9848 10310 15267 10362
rect 15319 10310 15331 10362
rect 15383 10310 15395 10362
rect 15447 10310 15459 10362
rect 15511 10310 15523 10362
rect 15575 10310 20994 10362
rect 21046 10310 21058 10362
rect 21110 10310 21122 10362
rect 21174 10310 21186 10362
rect 21238 10310 21250 10362
rect 21302 10310 24012 10362
rect 1104 10288 24012 10310
rect 13538 10208 13544 10260
rect 13596 10248 13602 10260
rect 18138 10248 18144 10260
rect 13596 10220 18144 10248
rect 13596 10208 13602 10220
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 20898 10208 20904 10260
rect 20956 10208 20962 10260
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 21450 10248 21456 10260
rect 21315 10220 21456 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 21450 10208 21456 10220
rect 21508 10208 21514 10260
rect 22002 10208 22008 10260
rect 22060 10208 22066 10260
rect 22094 10208 22100 10260
rect 22152 10208 22158 10260
rect 23477 10251 23535 10257
rect 23477 10217 23489 10251
rect 23523 10248 23535 10251
rect 24044 10248 24072 10628
rect 23523 10220 24072 10248
rect 23523 10217 23535 10220
rect 23477 10211 23535 10217
rect 8570 10180 8576 10192
rect 6932 10152 8576 10180
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5132 10084 5457 10112
rect 5132 10072 5138 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 6932 10112 6960 10152
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 14274 10140 14280 10192
rect 14332 10180 14338 10192
rect 20254 10180 20260 10192
rect 14332 10152 20260 10180
rect 14332 10140 14338 10152
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 20916 10180 20944 10208
rect 20916 10152 21128 10180
rect 6871 10084 6960 10112
rect 8113 10115 8171 10121
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 8113 10081 8125 10115
rect 8159 10112 8171 10115
rect 8202 10112 8208 10124
rect 8159 10084 8208 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 15838 10072 15844 10124
rect 15896 10072 15902 10124
rect 16025 10115 16083 10121
rect 16025 10081 16037 10115
rect 16071 10112 16083 10115
rect 16390 10112 16396 10124
rect 16071 10084 16396 10112
rect 16071 10081 16083 10084
rect 16025 10075 16083 10081
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 18506 10072 18512 10124
rect 18564 10112 18570 10124
rect 19242 10112 19248 10124
rect 18564 10084 19248 10112
rect 18564 10072 18570 10084
rect 19242 10072 19248 10084
rect 19300 10112 19306 10124
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 19300 10084 19809 10112
rect 19300 10072 19306 10084
rect 19797 10081 19809 10084
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 19978 10072 19984 10124
rect 20036 10112 20042 10124
rect 20533 10115 20591 10121
rect 20533 10112 20545 10115
rect 20036 10084 20545 10112
rect 20036 10072 20042 10084
rect 20533 10081 20545 10084
rect 20579 10081 20591 10115
rect 20533 10075 20591 10081
rect 20625 10115 20683 10121
rect 20625 10081 20637 10115
rect 20671 10081 20683 10115
rect 20625 10075 20683 10081
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 1627 10016 2774 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 2746 9976 2774 10016
rect 5258 10004 5264 10056
rect 5316 10004 5322 10056
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10044 5411 10047
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5399 10016 5733 10044
rect 5399 10013 5411 10016
rect 5353 10007 5411 10013
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10044 7067 10047
rect 7374 10044 7380 10056
rect 7055 10016 7380 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7834 10004 7840 10056
rect 7892 10004 7898 10056
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 7975 10016 8309 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8297 10007 8355 10013
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10044 15807 10047
rect 16114 10044 16120 10056
rect 15795 10016 16120 10044
rect 15795 10013 15807 10016
rect 15749 10007 15807 10013
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 17678 10004 17684 10056
rect 17736 10004 17742 10056
rect 19610 10004 19616 10056
rect 19668 10004 19674 10056
rect 20438 10004 20444 10056
rect 20496 10004 20502 10056
rect 6917 9979 6975 9985
rect 2746 9948 5028 9976
rect 1394 9868 1400 9920
rect 1452 9868 1458 9920
rect 4890 9868 4896 9920
rect 4948 9868 4954 9920
rect 5000 9908 5028 9948
rect 6917 9945 6929 9979
rect 6963 9976 6975 9979
rect 6963 9948 7512 9976
rect 6963 9945 6975 9948
rect 6917 9939 6975 9945
rect 7282 9908 7288 9920
rect 5000 9880 7288 9908
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 7374 9868 7380 9920
rect 7432 9868 7438 9920
rect 7484 9917 7512 9948
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 20640 9976 20668 10075
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 21100 10121 21128 10152
rect 22186 10140 22192 10192
rect 22244 10180 22250 10192
rect 22244 10152 23152 10180
rect 22244 10140 22250 10152
rect 23124 10124 23152 10152
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20772 10084 20913 10112
rect 20772 10072 20778 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 20901 10075 20959 10081
rect 21085 10115 21143 10121
rect 21085 10081 21097 10115
rect 21131 10081 21143 10115
rect 22465 10115 22523 10121
rect 22465 10112 22477 10115
rect 21085 10075 21143 10081
rect 21652 10084 22477 10112
rect 21652 10056 21680 10084
rect 22465 10081 22477 10084
rect 22511 10112 22523 10115
rect 22646 10112 22652 10124
rect 22511 10084 22652 10112
rect 22511 10081 22523 10084
rect 22465 10075 22523 10081
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 23014 10072 23020 10124
rect 23072 10072 23078 10124
rect 23106 10072 23112 10124
rect 23164 10072 23170 10124
rect 21634 10004 21640 10056
rect 21692 10004 21698 10056
rect 22281 10047 22339 10053
rect 22281 10044 22293 10047
rect 22066 10016 22293 10044
rect 19392 9948 20668 9976
rect 19392 9936 19398 9948
rect 21542 9936 21548 9988
rect 21600 9976 21606 9988
rect 21821 9979 21879 9985
rect 21821 9976 21833 9979
rect 21600 9948 21833 9976
rect 21600 9936 21606 9948
rect 21821 9945 21833 9948
rect 21867 9976 21879 9979
rect 22066 9976 22094 10016
rect 22281 10013 22293 10016
rect 22327 10044 22339 10047
rect 22327 10016 22600 10044
rect 22327 10013 22339 10016
rect 22281 10007 22339 10013
rect 21867 9948 22094 9976
rect 21867 9945 21879 9948
rect 21821 9939 21879 9945
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9877 7527 9911
rect 7469 9871 7527 9877
rect 15378 9868 15384 9920
rect 15436 9868 15442 9920
rect 17862 9868 17868 9920
rect 17920 9868 17926 9920
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 22572 9917 22600 10016
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 19245 9911 19303 9917
rect 19245 9908 19257 9911
rect 18012 9880 19257 9908
rect 18012 9868 18018 9880
rect 19245 9877 19257 9880
rect 19291 9877 19303 9911
rect 19245 9871 19303 9877
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9908 19763 9911
rect 20073 9911 20131 9917
rect 20073 9908 20085 9911
rect 19751 9880 20085 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 20073 9877 20085 9880
rect 20119 9877 20131 9911
rect 20073 9871 20131 9877
rect 22557 9911 22615 9917
rect 22557 9877 22569 9911
rect 22603 9877 22615 9911
rect 22557 9871 22615 9877
rect 22925 9911 22983 9917
rect 22925 9877 22937 9911
rect 22971 9908 22983 9911
rect 23290 9908 23296 9920
rect 22971 9880 23296 9908
rect 22971 9877 22983 9880
rect 22925 9871 22983 9877
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 1104 9818 24012 9840
rect 1104 9766 4473 9818
rect 4525 9766 4537 9818
rect 4589 9766 4601 9818
rect 4653 9766 4665 9818
rect 4717 9766 4729 9818
rect 4781 9766 10200 9818
rect 10252 9766 10264 9818
rect 10316 9766 10328 9818
rect 10380 9766 10392 9818
rect 10444 9766 10456 9818
rect 10508 9766 15927 9818
rect 15979 9766 15991 9818
rect 16043 9766 16055 9818
rect 16107 9766 16119 9818
rect 16171 9766 16183 9818
rect 16235 9766 21654 9818
rect 21706 9766 21718 9818
rect 21770 9766 21782 9818
rect 21834 9766 21846 9818
rect 21898 9766 21910 9818
rect 21962 9766 24012 9818
rect 1104 9744 24012 9766
rect 4890 9664 4896 9716
rect 4948 9664 4954 9716
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 7469 9707 7527 9713
rect 7469 9704 7481 9707
rect 7340 9676 7481 9704
rect 7340 9664 7346 9676
rect 7469 9673 7481 9676
rect 7515 9673 7527 9707
rect 7469 9667 7527 9673
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15657 9707 15715 9713
rect 15657 9704 15669 9707
rect 15436 9676 15669 9704
rect 15436 9664 15442 9676
rect 15657 9673 15669 9676
rect 15703 9673 15715 9707
rect 15657 9667 15715 9673
rect 17313 9707 17371 9713
rect 17313 9673 17325 9707
rect 17359 9673 17371 9707
rect 17313 9667 17371 9673
rect 4982 9596 4988 9648
rect 5040 9596 5046 9648
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7374 9636 7380 9648
rect 7055 9608 7380 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 13722 9636 13728 9648
rect 9876 9608 13728 9636
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 7392 9568 7420 9596
rect 7653 9571 7711 9577
rect 7653 9568 7665 9571
rect 7392 9540 7665 9568
rect 5629 9531 5687 9537
rect 7653 9537 7665 9540
rect 7699 9537 7711 9571
rect 9876 9568 9904 9608
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 17328 9636 17356 9667
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 23566 9704 23572 9716
rect 17920 9676 23572 9704
rect 17920 9664 17926 9676
rect 23566 9664 23572 9676
rect 23624 9664 23630 9716
rect 13872 9608 17356 9636
rect 17589 9639 17647 9645
rect 13872 9596 13878 9608
rect 17589 9605 17601 9639
rect 17635 9636 17647 9639
rect 17678 9636 17684 9648
rect 17635 9608 17684 9636
rect 17635 9605 17647 9608
rect 17589 9599 17647 9605
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 7653 9531 7711 9537
rect 9692 9540 9904 9568
rect 9968 9540 10425 9568
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9500 4859 9503
rect 4982 9500 4988 9512
rect 4847 9472 4988 9500
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5644 9500 5672 9531
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 5368 9472 7205 9500
rect 5368 9441 5396 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 8018 9500 8024 9512
rect 7423 9472 8024 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 5353 9435 5411 9441
rect 5353 9401 5365 9435
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 7009 9435 7067 9441
rect 7009 9401 7021 9435
rect 7055 9432 7067 9435
rect 9692 9432 9720 9540
rect 9968 9509 9996 9540
rect 10413 9537 10425 9540
rect 10459 9568 10471 9571
rect 10594 9568 10600 9580
rect 10459 9540 10600 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 10990 9571 11048 9577
rect 10990 9568 11002 9571
rect 10836 9540 11002 9568
rect 10836 9528 10842 9540
rect 10990 9537 11002 9540
rect 11036 9537 11048 9571
rect 10990 9531 11048 9537
rect 13446 9528 13452 9580
rect 13504 9528 13510 9580
rect 16574 9568 16580 9580
rect 15488 9540 16580 9568
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9500 10563 9503
rect 10686 9500 10692 9512
rect 10551 9472 10692 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 7055 9404 9720 9432
rect 9784 9432 9812 9463
rect 10520 9432 10548 9463
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 13265 9503 13323 9509
rect 13265 9500 13277 9503
rect 10928 9472 13277 9500
rect 10928 9460 10934 9472
rect 13265 9469 13277 9472
rect 13311 9469 13323 9503
rect 13265 9463 13323 9469
rect 9784 9404 10548 9432
rect 10781 9435 10839 9441
rect 7055 9401 7067 9404
rect 7009 9395 7067 9401
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 11238 9432 11244 9444
rect 10827 9404 11244 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 13280 9432 13308 9463
rect 13354 9460 13360 9512
rect 13412 9460 13418 9512
rect 15488 9509 15516 9540
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 16669 9571 16727 9577
rect 16669 9537 16681 9571
rect 16715 9568 16727 9571
rect 17221 9571 17279 9577
rect 17221 9568 17233 9571
rect 16715 9540 17233 9568
rect 16715 9537 16727 9540
rect 16669 9531 16727 9537
rect 17221 9537 17233 9540
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9568 17555 9571
rect 17954 9568 17960 9580
rect 17543 9540 17960 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 13740 9472 15485 9500
rect 13740 9432 13768 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15746 9500 15752 9512
rect 15611 9472 15752 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 13280 9404 13768 9432
rect 13817 9435 13875 9441
rect 13817 9401 13829 9435
rect 13863 9432 13875 9435
rect 16684 9432 16712 9531
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 23477 9571 23535 9577
rect 23477 9568 23489 9571
rect 22066 9540 23489 9568
rect 13863 9404 16712 9432
rect 18141 9435 18199 9441
rect 13863 9401 13875 9404
rect 13817 9395 13875 9401
rect 18141 9401 18153 9435
rect 18187 9432 18199 9435
rect 22066 9432 22094 9540
rect 23477 9537 23489 9540
rect 23523 9537 23535 9571
rect 23477 9531 23535 9537
rect 18187 9404 22094 9432
rect 18187 9401 18199 9404
rect 18141 9395 18199 9401
rect 23658 9392 23664 9444
rect 23716 9392 23722 9444
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 4856 9336 5457 9364
rect 4856 9324 4862 9336
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 7374 9364 7380 9376
rect 7331 9336 7380 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 9398 9324 9404 9376
rect 9456 9364 9462 9376
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 9456 9336 9597 9364
rect 9456 9324 9462 9336
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 10870 9324 10876 9376
rect 10928 9373 10934 9376
rect 10928 9367 10977 9373
rect 10928 9333 10931 9367
rect 10965 9333 10977 9367
rect 10928 9327 10977 9333
rect 10928 9324 10934 9327
rect 13906 9324 13912 9376
rect 13964 9324 13970 9376
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 16025 9367 16083 9373
rect 16025 9364 16037 9367
rect 15712 9336 16037 9364
rect 15712 9324 15718 9336
rect 16025 9333 16037 9336
rect 16071 9333 16083 9367
rect 16025 9327 16083 9333
rect 16206 9324 16212 9376
rect 16264 9324 16270 9376
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 17402 9324 17408 9376
rect 17460 9324 17466 9376
rect 1104 9274 24012 9296
rect 1104 9222 3813 9274
rect 3865 9222 3877 9274
rect 3929 9222 3941 9274
rect 3993 9222 4005 9274
rect 4057 9222 4069 9274
rect 4121 9222 9540 9274
rect 9592 9222 9604 9274
rect 9656 9222 9668 9274
rect 9720 9222 9732 9274
rect 9784 9222 9796 9274
rect 9848 9222 15267 9274
rect 15319 9222 15331 9274
rect 15383 9222 15395 9274
rect 15447 9222 15459 9274
rect 15511 9222 15523 9274
rect 15575 9222 20994 9274
rect 21046 9222 21058 9274
rect 21110 9222 21122 9274
rect 21174 9222 21186 9274
rect 21238 9222 21250 9274
rect 21302 9222 24012 9274
rect 1104 9200 24012 9222
rect 8018 9120 8024 9172
rect 8076 9120 8082 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 10962 9160 10968 9172
rect 8628 9132 10968 9160
rect 8628 9120 8634 9132
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 13412 9132 13737 9160
rect 13412 9120 13418 9132
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 15746 9120 15752 9172
rect 15804 9120 15810 9172
rect 842 9052 848 9104
rect 900 9092 906 9104
rect 1397 9095 1455 9101
rect 1397 9092 1409 9095
rect 900 9064 1409 9092
rect 900 9052 906 9064
rect 1397 9061 1409 9064
rect 1443 9061 1455 9095
rect 7745 9095 7803 9101
rect 7745 9092 7757 9095
rect 1397 9055 1455 9061
rect 6886 9064 7757 9092
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 6886 8956 6914 9064
rect 7745 9061 7757 9064
rect 7791 9061 7803 9095
rect 7745 9055 7803 9061
rect 1627 8928 6914 8956
rect 7929 8959 7987 8965
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8036 8956 8064 9120
rect 11609 9095 11667 9101
rect 11609 9092 11621 9095
rect 8496 9064 11621 9092
rect 8496 9033 8524 9064
rect 11609 9061 11621 9064
rect 11655 9061 11667 9095
rect 12802 9092 12808 9104
rect 11609 9055 11667 9061
rect 11992 9064 12808 9092
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 8481 8987 8539 8993
rect 8570 8984 8576 9036
rect 8628 8984 8634 9036
rect 9769 9027 9827 9033
rect 9769 8993 9781 9027
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 9024 11115 9027
rect 11992 9024 12020 9064
rect 12802 9052 12808 9064
rect 12860 9092 12866 9104
rect 14642 9092 14648 9104
rect 12860 9064 14648 9092
rect 12860 9052 12866 9064
rect 14642 9052 14648 9064
rect 14700 9052 14706 9104
rect 17773 9095 17831 9101
rect 17773 9061 17785 9095
rect 17819 9092 17831 9095
rect 17819 9064 22094 9092
rect 17819 9061 17831 9064
rect 17773 9055 17831 9061
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 11103 8996 12020 9024
rect 12084 8996 12173 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 7975 8928 8064 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9456 8928 9505 8956
rect 9456 8916 9462 8928
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9784 8956 9812 8987
rect 9784 8928 11100 8956
rect 9493 8919 9551 8925
rect 8389 8891 8447 8897
rect 8389 8857 8401 8891
rect 8435 8888 8447 8891
rect 10137 8891 10195 8897
rect 8435 8860 9168 8888
rect 8435 8857 8447 8860
rect 8389 8851 8447 8857
rect 9140 8829 9168 8860
rect 10137 8857 10149 8891
rect 10183 8857 10195 8891
rect 10137 8851 10195 8857
rect 10321 8891 10379 8897
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 10594 8888 10600 8900
rect 10367 8860 10600 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 9585 8823 9643 8829
rect 9585 8789 9597 8823
rect 9631 8820 9643 8823
rect 9953 8823 10011 8829
rect 9953 8820 9965 8823
rect 9631 8792 9965 8820
rect 9631 8789 9643 8792
rect 9585 8783 9643 8789
rect 9953 8789 9965 8792
rect 9999 8789 10011 8823
rect 10152 8820 10180 8851
rect 10594 8848 10600 8860
rect 10652 8848 10658 8900
rect 10781 8891 10839 8897
rect 10781 8857 10793 8891
rect 10827 8888 10839 8891
rect 10962 8888 10968 8900
rect 10827 8860 10968 8888
rect 10827 8857 10839 8860
rect 10781 8851 10839 8857
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 11072 8888 11100 8928
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11358 8959 11416 8965
rect 11358 8956 11370 8959
rect 11204 8928 11370 8956
rect 11204 8916 11210 8928
rect 11358 8925 11370 8928
rect 11404 8925 11416 8959
rect 11358 8919 11416 8925
rect 12084 8888 12112 8996
rect 12161 8993 12173 8996
rect 12207 9024 12219 9027
rect 13173 9027 13231 9033
rect 13173 9024 13185 9027
rect 12207 8996 13185 9024
rect 12207 8993 12219 8996
rect 12161 8987 12219 8993
rect 13173 8993 13185 8996
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 13906 9024 13912 9036
rect 13311 8996 13912 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 13188 8956 13216 8987
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 16206 8984 16212 9036
rect 16264 8984 16270 9036
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 19242 9024 19248 9036
rect 16448 8996 19248 9024
rect 16448 8984 16454 8996
rect 19242 8984 19248 8996
rect 19300 8984 19306 9036
rect 13722 8956 13728 8968
rect 13188 8928 13728 8956
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 17589 8959 17647 8965
rect 17589 8956 17601 8959
rect 17460 8928 17601 8956
rect 17460 8916 17466 8928
rect 17589 8925 17601 8928
rect 17635 8925 17647 8959
rect 22066 8956 22094 9064
rect 23477 8959 23535 8965
rect 23477 8956 23489 8959
rect 22066 8928 23489 8956
rect 17589 8919 17647 8925
rect 23477 8925 23489 8928
rect 23523 8925 23535 8959
rect 23477 8919 23535 8925
rect 11072 8860 12112 8888
rect 16117 8891 16175 8897
rect 16117 8857 16129 8891
rect 16163 8888 16175 8891
rect 16298 8888 16304 8900
rect 16163 8860 16304 8888
rect 16163 8857 16175 8860
rect 16117 8851 16175 8857
rect 16298 8848 16304 8860
rect 16356 8848 16362 8900
rect 10413 8823 10471 8829
rect 10413 8820 10425 8823
rect 10152 8792 10425 8820
rect 9953 8783 10011 8789
rect 10413 8789 10425 8792
rect 10459 8820 10471 8823
rect 10686 8820 10692 8832
rect 10459 8792 10692 8820
rect 10459 8789 10471 8792
rect 10413 8783 10471 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 11287 8823 11345 8829
rect 11287 8820 11299 8823
rect 10919 8792 11299 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 11287 8789 11299 8792
rect 11333 8789 11345 8823
rect 11287 8783 11345 8789
rect 11974 8780 11980 8832
rect 12032 8780 12038 8832
rect 12069 8823 12127 8829
rect 12069 8789 12081 8823
rect 12115 8820 12127 8823
rect 13354 8820 13360 8832
rect 12115 8792 13360 8820
rect 12115 8789 12127 8792
rect 12069 8783 12127 8789
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 23658 8780 23664 8832
rect 23716 8780 23722 8832
rect 1104 8730 24012 8752
rect 1104 8678 4473 8730
rect 4525 8678 4537 8730
rect 4589 8678 4601 8730
rect 4653 8678 4665 8730
rect 4717 8678 4729 8730
rect 4781 8678 10200 8730
rect 10252 8678 10264 8730
rect 10316 8678 10328 8730
rect 10380 8678 10392 8730
rect 10444 8678 10456 8730
rect 10508 8678 15927 8730
rect 15979 8678 15991 8730
rect 16043 8678 16055 8730
rect 16107 8678 16119 8730
rect 16171 8678 16183 8730
rect 16235 8678 21654 8730
rect 21706 8678 21718 8730
rect 21770 8678 21782 8730
rect 21834 8678 21846 8730
rect 21898 8678 21910 8730
rect 21962 8678 24012 8730
rect 1104 8656 24012 8678
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 5442 8616 5448 8628
rect 5307 8588 5448 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10870 8616 10876 8628
rect 10827 8588 10876 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 13446 8616 13452 8628
rect 13219 8588 13452 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 17460 8588 17877 8616
rect 17460 8576 17466 8588
rect 17865 8585 17877 8588
rect 17911 8585 17923 8619
rect 17865 8579 17923 8585
rect 18325 8619 18383 8625
rect 18325 8585 18337 8619
rect 18371 8616 18383 8619
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 18371 8588 18705 8616
rect 18371 8585 18383 8588
rect 18325 8579 18383 8585
rect 18693 8585 18705 8588
rect 18739 8585 18751 8619
rect 18693 8579 18751 8585
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 16908 8520 23520 8548
rect 16908 8508 16914 8520
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8480 4767 8483
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4755 8452 4905 8480
rect 4755 8449 4767 8452
rect 4709 8443 4767 8449
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5626 8480 5632 8492
rect 5123 8452 5632 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 10042 8440 10048 8492
rect 10100 8440 10106 8492
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 10778 8480 10784 8492
rect 10735 8452 10784 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11296 8452 11713 8480
rect 11296 8440 11302 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 13906 8480 13912 8492
rect 13587 8452 13912 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 15654 8480 15660 8492
rect 15611 8452 15660 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 16666 8440 16672 8492
rect 16724 8440 16730 8492
rect 18230 8440 18236 8492
rect 18288 8440 18294 8492
rect 19058 8440 19064 8492
rect 19116 8440 19122 8492
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8480 19211 8483
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 19199 8452 19533 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 19521 8449 19533 8452
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8480 22247 8483
rect 22554 8480 22560 8492
rect 22235 8452 22560 8480
rect 22235 8449 22247 8452
rect 22189 8443 22247 8449
rect 4522 8372 4528 8424
rect 4580 8372 4586 8424
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8381 11023 8415
rect 10965 8375 11023 8381
rect 4338 8304 4344 8356
rect 4396 8304 4402 8356
rect 9861 8347 9919 8353
rect 9861 8313 9873 8347
rect 9907 8344 9919 8347
rect 10594 8344 10600 8356
rect 9907 8316 10600 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 10594 8304 10600 8316
rect 10652 8304 10658 8356
rect 10980 8344 11008 8375
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 11204 8384 11621 8412
rect 11204 8372 11210 8384
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 11974 8372 11980 8424
rect 12032 8412 12038 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 12032 8384 12081 8412
rect 12032 8372 12038 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 13630 8372 13636 8424
rect 13688 8372 13694 8424
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 16390 8412 16396 8424
rect 13780 8384 16396 8412
rect 13780 8372 13786 8384
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 18506 8372 18512 8424
rect 18564 8372 18570 8424
rect 19242 8372 19248 8424
rect 19300 8372 19306 8424
rect 22020 8412 22048 8443
rect 22554 8440 22560 8452
rect 22612 8480 22618 8492
rect 22612 8452 22692 8480
rect 22612 8440 22618 8452
rect 22462 8412 22468 8424
rect 22020 8384 22468 8412
rect 22462 8372 22468 8384
rect 22520 8372 22526 8424
rect 22664 8421 22692 8452
rect 22922 8440 22928 8492
rect 22980 8489 22986 8492
rect 23492 8489 23520 8520
rect 22980 8483 23008 8489
rect 22996 8449 23008 8483
rect 22980 8443 23008 8449
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8449 23535 8483
rect 23477 8443 23535 8449
rect 22980 8440 22986 8443
rect 22649 8415 22707 8421
rect 22649 8381 22661 8415
rect 22695 8381 22707 8415
rect 22649 8375 22707 8381
rect 12342 8344 12348 8356
rect 10980 8316 12348 8344
rect 12342 8304 12348 8316
rect 12400 8304 12406 8356
rect 15749 8347 15807 8353
rect 15749 8313 15761 8347
rect 15795 8344 15807 8347
rect 17954 8344 17960 8356
rect 15795 8316 17960 8344
rect 15795 8313 15807 8316
rect 15749 8307 15807 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 20714 8344 20720 8356
rect 18064 8316 20720 8344
rect 4246 8236 4252 8288
rect 4304 8276 4310 8288
rect 5166 8276 5172 8288
rect 4304 8248 5172 8276
rect 4304 8236 4310 8248
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 10321 8279 10379 8285
rect 10321 8245 10333 8279
rect 10367 8276 10379 8279
rect 10502 8276 10508 8288
rect 10367 8248 10508 8276
rect 10367 8245 10379 8248
rect 10321 8239 10379 8245
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 16853 8279 16911 8285
rect 16853 8245 16865 8279
rect 16899 8276 16911 8279
rect 18064 8276 18092 8316
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 23661 8347 23719 8353
rect 23661 8344 23673 8347
rect 23440 8316 23673 8344
rect 23440 8304 23446 8316
rect 23661 8313 23673 8316
rect 23707 8313 23719 8347
rect 23661 8307 23719 8313
rect 16899 8248 18092 8276
rect 16899 8245 16911 8248
rect 16853 8239 16911 8245
rect 20898 8236 20904 8288
rect 20956 8236 20962 8288
rect 21726 8236 21732 8288
rect 21784 8276 21790 8288
rect 21821 8279 21879 8285
rect 21821 8276 21833 8279
rect 21784 8248 21833 8276
rect 21784 8236 21790 8248
rect 21821 8245 21833 8248
rect 21867 8245 21879 8279
rect 21821 8239 21879 8245
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 22281 8279 22339 8285
rect 22281 8276 22293 8279
rect 22244 8248 22293 8276
rect 22244 8236 22250 8248
rect 22281 8245 22293 8248
rect 22327 8245 22339 8279
rect 22281 8239 22339 8245
rect 22879 8279 22937 8285
rect 22879 8245 22891 8279
rect 22925 8276 22937 8279
rect 23014 8276 23020 8288
rect 22925 8248 23020 8276
rect 22925 8245 22937 8248
rect 22879 8239 22937 8245
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 1104 8186 24012 8208
rect 1104 8134 3813 8186
rect 3865 8134 3877 8186
rect 3929 8134 3941 8186
rect 3993 8134 4005 8186
rect 4057 8134 4069 8186
rect 4121 8134 9540 8186
rect 9592 8134 9604 8186
rect 9656 8134 9668 8186
rect 9720 8134 9732 8186
rect 9784 8134 9796 8186
rect 9848 8134 15267 8186
rect 15319 8134 15331 8186
rect 15383 8134 15395 8186
rect 15447 8134 15459 8186
rect 15511 8134 15523 8186
rect 15575 8134 20994 8186
rect 21046 8134 21058 8186
rect 21110 8134 21122 8186
rect 21174 8134 21186 8186
rect 21238 8134 21250 8186
rect 21302 8134 24012 8186
rect 1104 8112 24012 8134
rect 5626 8032 5632 8084
rect 5684 8032 5690 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 10226 8072 10232 8084
rect 10183 8044 10232 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 13449 8075 13507 8081
rect 13449 8041 13461 8075
rect 13495 8072 13507 8075
rect 13630 8072 13636 8084
rect 13495 8044 13636 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 13906 8032 13912 8084
rect 13964 8032 13970 8084
rect 15381 8075 15439 8081
rect 15381 8041 15393 8075
rect 15427 8072 15439 8075
rect 15838 8072 15844 8084
rect 15427 8044 15844 8072
rect 15427 8041 15439 8044
rect 15381 8035 15439 8041
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 19521 8075 19579 8081
rect 19521 8072 19533 8075
rect 16724 8044 19533 8072
rect 16724 8032 16730 8044
rect 19521 8041 19533 8044
rect 19567 8041 19579 8075
rect 19521 8035 19579 8041
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 22462 8072 22468 8084
rect 22152 8044 22468 8072
rect 22152 8032 22158 8044
rect 22462 8032 22468 8044
rect 22520 8072 22526 8084
rect 22557 8075 22615 8081
rect 22557 8072 22569 8075
rect 22520 8044 22569 8072
rect 22520 8032 22526 8044
rect 22557 8041 22569 8044
rect 22603 8041 22615 8075
rect 22557 8035 22615 8041
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 10873 8007 10931 8013
rect 10873 8004 10885 8007
rect 10100 7976 10885 8004
rect 10100 7964 10106 7976
rect 10873 7973 10885 7976
rect 10919 7973 10931 8007
rect 10873 7967 10931 7973
rect 15654 7964 15660 8016
rect 15712 8004 15718 8016
rect 15712 7976 15792 8004
rect 15712 7964 15718 7976
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4522 7936 4528 7948
rect 4479 7908 4528 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 4338 7828 4344 7880
rect 4396 7828 4402 7880
rect 4724 7868 4752 7899
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 4985 7939 5043 7945
rect 4985 7936 4997 7939
rect 4948 7908 4997 7936
rect 4948 7896 4954 7908
rect 4985 7905 4997 7908
rect 5031 7936 5043 7939
rect 5074 7936 5080 7948
rect 5031 7908 5080 7936
rect 5031 7905 5043 7908
rect 4985 7899 5043 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5350 7896 5356 7948
rect 5408 7936 5414 7948
rect 5997 7939 6055 7945
rect 5997 7936 6009 7939
rect 5408 7908 6009 7936
rect 5408 7896 5414 7908
rect 5997 7905 6009 7908
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 10502 7896 10508 7948
rect 10560 7896 10566 7948
rect 11057 7939 11115 7945
rect 11057 7905 11069 7939
rect 11103 7936 11115 7939
rect 11146 7936 11152 7948
rect 11103 7908 11152 7936
rect 11103 7905 11115 7908
rect 11057 7899 11115 7905
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 11238 7896 11244 7948
rect 11296 7896 11302 7948
rect 13538 7936 13544 7948
rect 13096 7908 13544 7936
rect 5718 7868 5724 7880
rect 4724 7840 5724 7868
rect 5718 7828 5724 7840
rect 5776 7868 5782 7880
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5776 7840 5825 7868
rect 5776 7828 5782 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7868 7251 7871
rect 7282 7868 7288 7880
rect 7239 7840 7288 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10686 7868 10692 7880
rect 10367 7840 10692 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 13096 7877 13124 7908
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 14642 7896 14648 7948
rect 14700 7896 14706 7948
rect 15562 7896 15568 7948
rect 15620 7896 15626 7948
rect 15764 7945 15792 7976
rect 21358 7964 21364 8016
rect 21416 8004 21422 8016
rect 21416 7976 22140 8004
rect 21416 7964 21422 7976
rect 15749 7939 15807 7945
rect 15749 7905 15761 7939
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 16942 7936 16948 7948
rect 16632 7908 16948 7936
rect 16632 7896 16638 7908
rect 16942 7896 16948 7908
rect 17000 7936 17006 7948
rect 20073 7939 20131 7945
rect 20073 7936 20085 7939
rect 17000 7908 20085 7936
rect 17000 7896 17006 7908
rect 20073 7905 20085 7908
rect 20119 7905 20131 7939
rect 20073 7899 20131 7905
rect 20898 7896 20904 7948
rect 20956 7896 20962 7948
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7936 21143 7939
rect 21131 7908 21588 7936
rect 21131 7905 21143 7908
rect 21085 7899 21143 7905
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7868 15715 7871
rect 16666 7868 16672 7880
rect 15703 7840 16672 7868
rect 15703 7837 15715 7840
rect 15657 7831 15715 7837
rect 7098 7800 7104 7812
rect 5552 7772 7104 7800
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2590 7732 2596 7744
rect 1627 7704 2596 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 5074 7692 5080 7744
rect 5132 7692 5138 7744
rect 5166 7692 5172 7744
rect 5224 7692 5230 7744
rect 5552 7741 5580 7772
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 13170 7760 13176 7812
rect 13228 7800 13234 7812
rect 13265 7803 13323 7809
rect 13265 7800 13277 7803
rect 13228 7772 13277 7800
rect 13228 7760 13234 7772
rect 13265 7769 13277 7772
rect 13311 7800 13323 7803
rect 13740 7800 13768 7831
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 21560 7812 21588 7908
rect 21726 7896 21732 7948
rect 21784 7896 21790 7948
rect 22112 7945 22140 7976
rect 21821 7939 21879 7945
rect 21821 7905 21833 7939
rect 21867 7905 21879 7939
rect 21821 7899 21879 7905
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7905 22155 7939
rect 22097 7899 22155 7905
rect 13311 7772 13768 7800
rect 13311 7769 13323 7772
rect 13265 7763 13323 7769
rect 5537 7735 5595 7741
rect 5537 7701 5549 7735
rect 5583 7701 5595 7735
rect 13740 7732 13768 7772
rect 14458 7760 14464 7812
rect 14516 7800 14522 7812
rect 14516 7772 15010 7800
rect 14516 7760 14522 7772
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13740 7704 14105 7732
rect 5537 7695 5595 7701
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 14550 7692 14556 7744
rect 14608 7692 14614 7744
rect 14982 7732 15010 7772
rect 15194 7760 15200 7812
rect 15252 7800 15258 7812
rect 15381 7803 15439 7809
rect 15381 7800 15393 7803
rect 15252 7772 15393 7800
rect 15252 7760 15258 7772
rect 15381 7769 15393 7772
rect 15427 7769 15439 7803
rect 15381 7763 15439 7769
rect 19889 7803 19947 7809
rect 19889 7769 19901 7803
rect 19935 7800 19947 7803
rect 19935 7772 21312 7800
rect 19935 7769 19947 7772
rect 19889 7763 19947 7769
rect 16482 7732 16488 7744
rect 14982 7704 16488 7732
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 19981 7735 20039 7741
rect 19981 7701 19993 7735
rect 20027 7732 20039 7735
rect 20441 7735 20499 7741
rect 20441 7732 20453 7735
rect 20027 7704 20453 7732
rect 20027 7701 20039 7704
rect 19981 7695 20039 7701
rect 20441 7701 20453 7704
rect 20487 7701 20499 7735
rect 20441 7695 20499 7701
rect 20809 7735 20867 7741
rect 20809 7701 20821 7735
rect 20855 7732 20867 7735
rect 21082 7732 21088 7744
rect 20855 7704 21088 7732
rect 20855 7701 20867 7704
rect 20809 7695 20867 7701
rect 21082 7692 21088 7704
rect 21140 7692 21146 7744
rect 21284 7741 21312 7772
rect 21542 7760 21548 7812
rect 21600 7800 21606 7812
rect 21836 7800 21864 7899
rect 23106 7896 23112 7948
rect 23164 7896 23170 7948
rect 22186 7868 22192 7880
rect 21600 7772 21864 7800
rect 21928 7840 22192 7868
rect 21600 7760 21606 7772
rect 21269 7735 21327 7741
rect 21269 7701 21281 7735
rect 21315 7701 21327 7735
rect 21269 7695 21327 7701
rect 21637 7735 21695 7741
rect 21637 7701 21649 7735
rect 21683 7732 21695 7735
rect 21928 7732 21956 7840
rect 22186 7828 22192 7840
rect 22244 7828 22250 7880
rect 22281 7871 22339 7877
rect 22281 7837 22293 7871
rect 22327 7837 22339 7871
rect 22281 7831 22339 7837
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7868 22983 7871
rect 23474 7868 23480 7880
rect 23532 7877 23538 7880
rect 23532 7871 23560 7877
rect 22971 7840 23480 7868
rect 22971 7837 22983 7840
rect 22925 7831 22983 7837
rect 22002 7760 22008 7812
rect 22060 7800 22066 7812
rect 22296 7800 22324 7831
rect 23474 7828 23480 7840
rect 23548 7837 23560 7871
rect 23532 7831 23560 7837
rect 23532 7828 23538 7831
rect 22060 7772 22324 7800
rect 22060 7760 22066 7772
rect 21683 7704 21956 7732
rect 21683 7701 21695 7704
rect 21637 7695 21695 7701
rect 22462 7692 22468 7744
rect 22520 7692 22526 7744
rect 23017 7735 23075 7741
rect 23017 7701 23029 7735
rect 23063 7732 23075 7735
rect 23431 7735 23489 7741
rect 23431 7732 23443 7735
rect 23063 7704 23443 7732
rect 23063 7701 23075 7704
rect 23017 7695 23075 7701
rect 23431 7701 23443 7704
rect 23477 7701 23489 7735
rect 23431 7695 23489 7701
rect 1104 7642 24012 7664
rect 1104 7590 4473 7642
rect 4525 7590 4537 7642
rect 4589 7590 4601 7642
rect 4653 7590 4665 7642
rect 4717 7590 4729 7642
rect 4781 7590 10200 7642
rect 10252 7590 10264 7642
rect 10316 7590 10328 7642
rect 10380 7590 10392 7642
rect 10444 7590 10456 7642
rect 10508 7590 15927 7642
rect 15979 7590 15991 7642
rect 16043 7590 16055 7642
rect 16107 7590 16119 7642
rect 16171 7590 16183 7642
rect 16235 7590 21654 7642
rect 21706 7590 21718 7642
rect 21770 7590 21782 7642
rect 21834 7590 21846 7642
rect 21898 7590 21910 7642
rect 21962 7590 24012 7642
rect 1104 7568 24012 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 3697 7531 3755 7537
rect 1627 7500 3464 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 2590 7420 2596 7472
rect 2648 7460 2654 7472
rect 3329 7463 3387 7469
rect 3329 7460 3341 7463
rect 2648 7432 3341 7460
rect 2648 7420 2654 7432
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 2700 7401 2728 7432
rect 3329 7429 3341 7432
rect 3375 7429 3387 7463
rect 3329 7423 3387 7429
rect 2700 7395 2778 7401
rect 2700 7364 2732 7395
rect 2720 7361 2732 7364
rect 2766 7361 2778 7395
rect 2720 7355 2778 7361
rect 2823 7395 2881 7401
rect 2823 7361 2835 7395
rect 2869 7392 2881 7395
rect 3237 7395 3295 7401
rect 3237 7392 3249 7395
rect 2869 7364 3249 7392
rect 2869 7361 2881 7364
rect 2823 7355 2881 7361
rect 3237 7361 3249 7364
rect 3283 7361 3295 7395
rect 3436 7392 3464 7500
rect 3697 7497 3709 7531
rect 3743 7528 3755 7531
rect 4338 7528 4344 7540
rect 3743 7500 4344 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 4338 7488 4344 7500
rect 4396 7528 4402 7540
rect 4396 7500 5028 7528
rect 4396 7488 4402 7500
rect 5000 7469 5028 7500
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 5132 7500 5365 7528
rect 5132 7488 5138 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 7282 7488 7288 7540
rect 7340 7488 7346 7540
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 13262 7528 13268 7540
rect 9079 7500 13268 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 14047 7531 14105 7537
rect 14047 7497 14059 7531
rect 14093 7528 14105 7531
rect 14550 7528 14556 7540
rect 14093 7500 14556 7528
rect 14093 7497 14105 7500
rect 14047 7491 14105 7497
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 22554 7488 22560 7540
rect 22612 7488 22618 7540
rect 22922 7488 22928 7540
rect 22980 7488 22986 7540
rect 23014 7488 23020 7540
rect 23072 7488 23078 7540
rect 23477 7531 23535 7537
rect 23477 7497 23489 7531
rect 23523 7497 23535 7531
rect 23477 7491 23535 7497
rect 4525 7463 4583 7469
rect 4525 7460 4537 7463
rect 3896 7432 4537 7460
rect 3896 7401 3924 7432
rect 4525 7429 4537 7432
rect 4571 7429 4583 7463
rect 4525 7423 4583 7429
rect 4985 7463 5043 7469
rect 4985 7429 4997 7463
rect 5031 7429 5043 7463
rect 4985 7423 5043 7429
rect 3896 7395 3974 7401
rect 3896 7392 3928 7395
rect 3436 7364 3928 7392
rect 3237 7355 3295 7361
rect 3916 7361 3928 7364
rect 3962 7361 3974 7395
rect 3916 7355 3974 7361
rect 4019 7395 4077 7401
rect 4019 7361 4031 7395
rect 4065 7392 4077 7395
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4065 7364 4445 7392
rect 4065 7361 4077 7364
rect 4019 7355 4077 7361
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 4433 7355 4491 7361
rect 4908 7364 5181 7392
rect 3145 7327 3203 7333
rect 3145 7293 3157 7327
rect 3191 7324 3203 7327
rect 3191 7296 4200 7324
rect 3191 7293 3203 7296
rect 3145 7287 3203 7293
rect 4172 7188 4200 7296
rect 4246 7284 4252 7336
rect 4304 7284 4310 7336
rect 4798 7216 4804 7268
rect 4856 7256 4862 7268
rect 4908 7265 4936 7364
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5350 7352 5356 7404
rect 5408 7392 5414 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5408 7364 5825 7392
rect 5408 7352 5414 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 5813 7355 5871 7361
rect 6196 7364 7205 7392
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 6196 7333 6224 7364
rect 7193 7361 7205 7364
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7524 7364 7849 7392
rect 7524 7352 7530 7364
rect 7837 7361 7849 7364
rect 7883 7392 7895 7395
rect 9125 7395 9183 7401
rect 7883 7364 8984 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7293 6239 7327
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 6181 7287 6239 7293
rect 6886 7296 7389 7324
rect 4893 7259 4951 7265
rect 4893 7256 4905 7259
rect 4856 7228 4905 7256
rect 4856 7216 4862 7228
rect 4893 7225 4905 7228
rect 4939 7225 4951 7259
rect 4893 7219 4951 7225
rect 5258 7216 5264 7268
rect 5316 7256 5322 7268
rect 6886 7256 6914 7296
rect 7377 7293 7389 7296
rect 7423 7324 7435 7327
rect 7926 7324 7932 7336
rect 7423 7296 7932 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 7926 7284 7932 7296
rect 7984 7324 7990 7336
rect 8202 7324 8208 7336
rect 7984 7296 8208 7324
rect 7984 7284 7990 7296
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8754 7284 8760 7336
rect 8812 7284 8818 7336
rect 8956 7333 8984 7364
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9306 7392 9312 7404
rect 9171 7364 9312 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9306 7352 9312 7364
rect 9364 7392 9370 7404
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9364 7364 9413 7392
rect 9364 7352 9370 7364
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 13976 7395 14034 7401
rect 13976 7361 13988 7395
rect 14022 7392 14034 7395
rect 14458 7392 14464 7404
rect 14022 7364 14464 7392
rect 14022 7361 14034 7364
rect 13976 7355 14034 7361
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 15289 7395 15347 7401
rect 15289 7392 15301 7395
rect 15252 7364 15301 7392
rect 15252 7352 15258 7364
rect 15289 7361 15301 7364
rect 15335 7361 15347 7395
rect 15289 7355 15347 7361
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15933 7395 15991 7401
rect 15933 7392 15945 7395
rect 15620 7364 15945 7392
rect 15620 7352 15626 7364
rect 15933 7361 15945 7364
rect 15979 7392 15991 7395
rect 16298 7392 16304 7404
rect 15979 7364 16304 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 18690 7352 18696 7404
rect 18748 7352 18754 7404
rect 21358 7352 21364 7404
rect 21416 7392 21422 7404
rect 21453 7395 21511 7401
rect 21453 7392 21465 7395
rect 21416 7364 21465 7392
rect 21416 7352 21422 7364
rect 21453 7361 21465 7364
rect 21499 7361 21511 7395
rect 21453 7355 21511 7361
rect 22186 7352 22192 7404
rect 22244 7392 22250 7404
rect 22572 7392 22600 7488
rect 22940 7460 22968 7488
rect 23492 7460 23520 7491
rect 22940 7432 23520 7460
rect 22244 7364 22600 7392
rect 22244 7352 22250 7364
rect 23658 7352 23664 7404
rect 23716 7352 23722 7404
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 18785 7327 18843 7333
rect 18785 7293 18797 7327
rect 18831 7324 18843 7327
rect 18874 7324 18880 7336
rect 18831 7296 18880 7324
rect 18831 7293 18843 7296
rect 18785 7287 18843 7293
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 19058 7284 19064 7336
rect 19116 7284 19122 7336
rect 21082 7284 21088 7336
rect 21140 7284 21146 7336
rect 21545 7327 21603 7333
rect 21545 7293 21557 7327
rect 21591 7324 21603 7327
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21591 7296 21833 7324
rect 21591 7293 21603 7296
rect 21545 7287 21603 7293
rect 21821 7293 21833 7296
rect 21867 7324 21879 7327
rect 22002 7324 22008 7336
rect 21867 7296 22008 7324
rect 21867 7293 21879 7296
rect 21821 7287 21879 7293
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 22094 7284 22100 7336
rect 22152 7284 22158 7336
rect 23198 7284 23204 7336
rect 23256 7284 23262 7336
rect 5316 7228 6914 7256
rect 15473 7259 15531 7265
rect 5316 7216 5322 7228
rect 15473 7225 15485 7259
rect 15519 7256 15531 7259
rect 16390 7256 16396 7268
rect 15519 7228 16396 7256
rect 15519 7225 15531 7228
rect 15473 7219 15531 7225
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 5442 7188 5448 7200
rect 4172 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 7006 7188 7012 7200
rect 6871 7160 7012 7188
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 8018 7148 8024 7200
rect 8076 7148 8082 7200
rect 8386 7148 8392 7200
rect 8444 7188 8450 7200
rect 8849 7191 8907 7197
rect 8849 7188 8861 7191
rect 8444 7160 8861 7188
rect 8444 7148 8450 7160
rect 8849 7157 8861 7160
rect 8895 7157 8907 7191
rect 8849 7151 8907 7157
rect 9217 7191 9275 7197
rect 9217 7157 9229 7191
rect 9263 7188 9275 7191
rect 9306 7188 9312 7200
rect 9263 7160 9312 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 16117 7191 16175 7197
rect 16117 7157 16129 7191
rect 16163 7188 16175 7191
rect 17034 7188 17040 7200
rect 16163 7160 17040 7188
rect 16163 7157 16175 7160
rect 16117 7151 16175 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 1104 7098 24012 7120
rect 1104 7046 3813 7098
rect 3865 7046 3877 7098
rect 3929 7046 3941 7098
rect 3993 7046 4005 7098
rect 4057 7046 4069 7098
rect 4121 7046 9540 7098
rect 9592 7046 9604 7098
rect 9656 7046 9668 7098
rect 9720 7046 9732 7098
rect 9784 7046 9796 7098
rect 9848 7046 15267 7098
rect 15319 7046 15331 7098
rect 15383 7046 15395 7098
rect 15447 7046 15459 7098
rect 15511 7046 15523 7098
rect 15575 7046 20994 7098
rect 21046 7046 21058 7098
rect 21110 7046 21122 7098
rect 21174 7046 21186 7098
rect 21238 7046 21250 7098
rect 21302 7046 24012 7098
rect 1104 7024 24012 7046
rect 4801 6987 4859 6993
rect 4801 6953 4813 6987
rect 4847 6984 4859 6987
rect 5166 6984 5172 6996
rect 4847 6956 5172 6984
rect 4847 6953 4859 6956
rect 4801 6947 4859 6953
rect 5166 6944 5172 6956
rect 5224 6944 5230 6996
rect 5258 6944 5264 6996
rect 5316 6984 5322 6996
rect 5442 6984 5448 6996
rect 5316 6956 5448 6984
rect 5316 6944 5322 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 7466 6944 7472 6996
rect 7524 6944 7530 6996
rect 16298 6944 16304 6996
rect 16356 6944 16362 6996
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 4433 6919 4491 6925
rect 4433 6916 4445 6919
rect 4396 6888 4445 6916
rect 4396 6876 4402 6888
rect 4433 6885 4445 6888
rect 4479 6885 4491 6919
rect 13538 6916 13544 6928
rect 4433 6879 4491 6885
rect 6932 6888 7144 6916
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 4798 6848 4804 6860
rect 4663 6820 4804 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 6932 6857 6960 6888
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 5040 6820 6929 6848
rect 5040 6808 5046 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 7116 6848 7144 6888
rect 12912 6888 13544 6916
rect 8570 6848 8576 6860
rect 7116 6820 8576 6848
rect 6917 6811 6975 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 7098 6740 7104 6792
rect 7156 6740 7162 6792
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7432 6752 7757 6780
rect 7432 6740 7438 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9582 6780 9588 6792
rect 8812 6752 9588 6780
rect 8812 6740 8818 6752
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 10962 6780 10968 6792
rect 10919 6752 10968 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 12912 6789 12940 6888
rect 13538 6876 13544 6888
rect 13596 6916 13602 6928
rect 13725 6919 13783 6925
rect 13725 6916 13737 6919
rect 13596 6888 13737 6916
rect 13596 6876 13602 6888
rect 13725 6885 13737 6888
rect 13771 6885 13783 6919
rect 18138 6916 18144 6928
rect 13725 6879 13783 6885
rect 17972 6888 18144 6916
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6749 12955 6783
rect 13004 6780 13032 6811
rect 13262 6808 13268 6860
rect 13320 6808 13326 6860
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6848 15715 6851
rect 16942 6848 16948 6860
rect 15703 6820 16948 6848
rect 15703 6817 15715 6820
rect 15657 6811 15715 6817
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6848 17831 6851
rect 17972 6848 18000 6888
rect 18138 6876 18144 6888
rect 18196 6916 18202 6928
rect 19242 6916 19248 6928
rect 18196 6888 19248 6916
rect 18196 6876 18202 6888
rect 19242 6876 19248 6888
rect 19300 6916 19306 6928
rect 21542 6916 21548 6928
rect 19300 6888 21548 6916
rect 19300 6876 19306 6888
rect 21542 6876 21548 6888
rect 21600 6876 21606 6928
rect 22186 6876 22192 6928
rect 22244 6876 22250 6928
rect 17819 6820 18000 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 19061 6851 19119 6857
rect 19061 6848 19073 6851
rect 18748 6820 19073 6848
rect 18748 6808 18754 6820
rect 19061 6817 19073 6820
rect 19107 6848 19119 6851
rect 21361 6851 21419 6857
rect 21361 6848 21373 6851
rect 19107 6820 21373 6848
rect 19107 6817 19119 6820
rect 19061 6811 19119 6817
rect 21361 6817 21373 6820
rect 21407 6817 21419 6851
rect 21361 6811 21419 6817
rect 22005 6851 22063 6857
rect 22005 6817 22017 6851
rect 22051 6848 22063 6851
rect 22094 6848 22100 6860
rect 22051 6820 22100 6848
rect 22051 6817 22063 6820
rect 22005 6811 22063 6817
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 13170 6780 13176 6792
rect 13004 6752 13176 6780
rect 12897 6743 12955 6749
rect 13170 6740 13176 6752
rect 13228 6780 13234 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13228 6752 13553 6780
rect 13228 6740 13234 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 17957 6783 18015 6789
rect 17957 6780 17969 6783
rect 17635 6752 17969 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 17957 6749 17969 6752
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 18874 6740 18880 6792
rect 18932 6740 18938 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 22462 6780 22468 6792
rect 21591 6752 22468 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6780 23535 6783
rect 23566 6780 23572 6792
rect 23523 6752 23572 6780
rect 23523 6749 23535 6752
rect 23477 6743 23535 6749
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 15381 6715 15439 6721
rect 15381 6681 15393 6715
rect 15427 6712 15439 6715
rect 15654 6712 15660 6724
rect 15427 6684 15660 6712
rect 15427 6681 15439 6684
rect 15381 6675 15439 6681
rect 15654 6672 15660 6684
rect 15712 6672 15718 6724
rect 21729 6715 21787 6721
rect 21729 6681 21741 6715
rect 21775 6712 21787 6715
rect 21821 6715 21879 6721
rect 21821 6712 21833 6715
rect 21775 6684 21833 6712
rect 21775 6681 21787 6684
rect 21729 6675 21787 6681
rect 21821 6681 21833 6684
rect 21867 6681 21879 6715
rect 21821 6675 21879 6681
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7561 6647 7619 6653
rect 7561 6644 7573 6647
rect 7064 6616 7573 6644
rect 7064 6604 7070 6616
rect 7561 6613 7573 6616
rect 7607 6613 7619 6647
rect 7561 6607 7619 6613
rect 8570 6604 8576 6656
rect 8628 6604 8634 6656
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 9950 6644 9956 6656
rect 9815 6616 9956 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6644 13415 6647
rect 13446 6644 13452 6656
rect 13403 6616 13452 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6644 15071 6647
rect 15194 6644 15200 6656
rect 15059 6616 15200 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15470 6604 15476 6656
rect 15528 6604 15534 6656
rect 16666 6604 16672 6656
rect 16724 6604 16730 6656
rect 16761 6647 16819 6653
rect 16761 6613 16773 6647
rect 16807 6644 16819 6647
rect 17129 6647 17187 6653
rect 17129 6644 17141 6647
rect 16807 6616 17141 6644
rect 16807 6613 16819 6616
rect 16761 6607 16819 6613
rect 17129 6613 17141 6616
rect 17175 6613 17187 6647
rect 17129 6607 17187 6613
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17497 6647 17555 6653
rect 17497 6644 17509 6647
rect 17276 6616 17509 6644
rect 17276 6604 17282 6616
rect 17497 6613 17509 6616
rect 17543 6613 17555 6647
rect 17497 6607 17555 6613
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 18693 6647 18751 6653
rect 18693 6644 18705 6647
rect 18564 6616 18705 6644
rect 18564 6604 18570 6616
rect 18693 6613 18705 6616
rect 18739 6613 18751 6647
rect 18693 6607 18751 6613
rect 23658 6604 23664 6656
rect 23716 6604 23722 6656
rect 1104 6554 24012 6576
rect 1104 6502 4473 6554
rect 4525 6502 4537 6554
rect 4589 6502 4601 6554
rect 4653 6502 4665 6554
rect 4717 6502 4729 6554
rect 4781 6502 10200 6554
rect 10252 6502 10264 6554
rect 10316 6502 10328 6554
rect 10380 6502 10392 6554
rect 10444 6502 10456 6554
rect 10508 6502 15927 6554
rect 15979 6502 15991 6554
rect 16043 6502 16055 6554
rect 16107 6502 16119 6554
rect 16171 6502 16183 6554
rect 16235 6502 21654 6554
rect 21706 6502 21718 6554
rect 21770 6502 21782 6554
rect 21834 6502 21846 6554
rect 21898 6502 21910 6554
rect 21962 6502 24012 6554
rect 1104 6480 24012 6502
rect 8113 6443 8171 6449
rect 8113 6409 8125 6443
rect 8159 6440 8171 6443
rect 8665 6443 8723 6449
rect 8665 6440 8677 6443
rect 8159 6412 8677 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 8665 6409 8677 6412
rect 8711 6409 8723 6443
rect 8665 6403 8723 6409
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 9640 6412 9689 6440
rect 9640 6400 9646 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 9677 6403 9735 6409
rect 10137 6443 10195 6449
rect 10137 6409 10149 6443
rect 10183 6440 10195 6443
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10183 6412 10517 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 10870 6440 10876 6452
rect 10744 6412 10876 6440
rect 10744 6400 10750 6412
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 10962 6400 10968 6452
rect 11020 6400 11026 6452
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13538 6440 13544 6452
rect 13219 6412 13544 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 15470 6440 15476 6452
rect 15427 6412 15476 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 18230 6400 18236 6452
rect 18288 6440 18294 6452
rect 18785 6443 18843 6449
rect 18785 6440 18797 6443
rect 18288 6412 18797 6440
rect 18288 6400 18294 6412
rect 18785 6409 18797 6412
rect 18831 6409 18843 6443
rect 18785 6403 18843 6409
rect 23474 6400 23480 6452
rect 23532 6400 23538 6452
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 12805 6375 12863 6381
rect 8812 6344 10272 6372
rect 8812 6332 8818 6344
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8478 6304 8484 6316
rect 8251 6276 8484 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8588 6276 9045 6304
rect 4982 6196 4988 6248
rect 5040 6236 5046 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 5040 6208 7941 6236
rect 5040 6196 5046 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 7929 6199 7987 6205
rect 8294 6196 8300 6248
rect 8352 6236 8358 6248
rect 8588 6236 8616 6276
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 8352 6208 8616 6236
rect 8352 6196 8358 6208
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 10244 6245 10272 6344
rect 12805 6341 12817 6375
rect 12851 6372 12863 6375
rect 14274 6372 14280 6384
rect 12851 6344 14280 6372
rect 12851 6341 12863 6344
rect 12805 6335 12863 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 18506 6332 18512 6384
rect 18564 6332 18570 6384
rect 19242 6332 19248 6384
rect 19300 6332 19306 6384
rect 10870 6264 10876 6316
rect 10928 6264 10934 6316
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6273 13691 6307
rect 13633 6267 13691 6273
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8720 6208 9137 6236
rect 8720 6196 8726 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9217 6239 9275 6245
rect 9217 6205 9229 6239
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 11057 6239 11115 6245
rect 11057 6236 11069 6239
rect 10229 6199 10287 6205
rect 10336 6208 11069 6236
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 8573 6171 8631 6177
rect 8573 6168 8585 6171
rect 8444 6140 8585 6168
rect 8444 6128 8450 6140
rect 8573 6137 8585 6140
rect 8619 6137 8631 6171
rect 9232 6168 9260 6199
rect 10336 6168 10364 6208
rect 11057 6205 11069 6208
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 12526 6196 12532 6248
rect 12584 6196 12590 6248
rect 12710 6196 12716 6248
rect 12768 6196 12774 6248
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 13541 6239 13599 6245
rect 13541 6236 13553 6239
rect 13320 6208 13553 6236
rect 13320 6196 13326 6208
rect 13541 6205 13553 6208
rect 13587 6205 13599 6239
rect 13648 6236 13676 6267
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13872 6276 14105 6304
rect 13872 6264 13878 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 15746 6264 15752 6316
rect 15804 6264 15810 6316
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6304 15899 6307
rect 16209 6307 16267 6313
rect 16209 6304 16221 6307
rect 15887 6276 16221 6304
rect 15887 6273 15899 6276
rect 15841 6267 15899 6273
rect 16209 6273 16221 6276
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 18966 6304 18972 6316
rect 18739 6276 18972 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19150 6264 19156 6316
rect 19208 6264 19214 6316
rect 19260 6304 19288 6332
rect 19260 6276 19380 6304
rect 14185 6239 14243 6245
rect 14185 6236 14197 6239
rect 13648 6208 14197 6236
rect 13541 6199 13599 6205
rect 14185 6205 14197 6208
rect 14231 6236 14243 6239
rect 14366 6236 14372 6248
rect 14231 6208 14372 6236
rect 14231 6205 14243 6208
rect 14185 6199 14243 6205
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 16025 6239 16083 6245
rect 16025 6205 16037 6239
rect 16071 6236 16083 6239
rect 18138 6236 18144 6248
rect 16071 6208 18144 6236
rect 16071 6205 16083 6208
rect 16025 6199 16083 6205
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 19242 6196 19248 6248
rect 19300 6196 19306 6248
rect 19352 6245 19380 6276
rect 19978 6264 19984 6316
rect 20036 6264 20042 6316
rect 23658 6264 23664 6316
rect 23716 6264 23722 6316
rect 19337 6239 19395 6245
rect 19337 6205 19349 6239
rect 19383 6205 19395 6239
rect 19337 6199 19395 6205
rect 20073 6239 20131 6245
rect 20073 6205 20085 6239
rect 20119 6236 20131 6239
rect 20162 6236 20168 6248
rect 20119 6208 20168 6236
rect 20119 6205 20131 6208
rect 20073 6199 20131 6205
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 8573 6131 8631 6137
rect 9140 6140 10364 6168
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 9140 6100 9168 6140
rect 18874 6128 18880 6180
rect 18932 6168 18938 6180
rect 19613 6171 19671 6177
rect 19613 6168 19625 6171
rect 18932 6140 19625 6168
rect 18932 6128 18938 6140
rect 19613 6137 19625 6140
rect 19659 6137 19671 6171
rect 19613 6131 19671 6137
rect 7984 6072 9168 6100
rect 13265 6103 13323 6109
rect 7984 6060 7990 6072
rect 13265 6069 13277 6103
rect 13311 6100 13323 6103
rect 13354 6100 13360 6112
rect 13311 6072 13360 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 14461 6103 14519 6109
rect 14461 6069 14473 6103
rect 14507 6100 14519 6103
rect 15838 6100 15844 6112
rect 14507 6072 15844 6100
rect 14507 6069 14519 6072
rect 14461 6063 14519 6069
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 17586 6060 17592 6112
rect 17644 6100 17650 6112
rect 18325 6103 18383 6109
rect 18325 6100 18337 6103
rect 17644 6072 18337 6100
rect 17644 6060 17650 6072
rect 18325 6069 18337 6072
rect 18371 6069 18383 6103
rect 18325 6063 18383 6069
rect 1104 6010 24012 6032
rect 1104 5958 3813 6010
rect 3865 5958 3877 6010
rect 3929 5958 3941 6010
rect 3993 5958 4005 6010
rect 4057 5958 4069 6010
rect 4121 5958 9540 6010
rect 9592 5958 9604 6010
rect 9656 5958 9668 6010
rect 9720 5958 9732 6010
rect 9784 5958 9796 6010
rect 9848 5958 15267 6010
rect 15319 5958 15331 6010
rect 15383 5958 15395 6010
rect 15447 5958 15459 6010
rect 15511 5958 15523 6010
rect 15575 5958 20994 6010
rect 21046 5958 21058 6010
rect 21110 5958 21122 6010
rect 21174 5958 21186 6010
rect 21238 5958 21250 6010
rect 21302 5958 24012 6010
rect 1104 5936 24012 5958
rect 5537 5899 5595 5905
rect 5537 5865 5549 5899
rect 5583 5896 5595 5899
rect 7374 5896 7380 5908
rect 5583 5868 7380 5896
rect 5583 5865 5595 5868
rect 5537 5859 5595 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 8662 5856 8668 5908
rect 8720 5856 8726 5908
rect 10870 5856 10876 5908
rect 10928 5896 10934 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 10928 5868 11069 5896
rect 10928 5856 10934 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 12710 5856 12716 5908
rect 12768 5905 12774 5908
rect 12768 5899 12817 5905
rect 12768 5865 12771 5899
rect 12805 5865 12817 5899
rect 12768 5859 12817 5865
rect 12768 5856 12774 5859
rect 17218 5856 17224 5908
rect 17276 5856 17282 5908
rect 18693 5899 18751 5905
rect 18693 5865 18705 5899
rect 18739 5896 18751 5899
rect 19150 5896 19156 5908
rect 18739 5868 19156 5896
rect 18739 5865 18751 5868
rect 18693 5859 18751 5865
rect 19150 5856 19156 5868
rect 19208 5856 19214 5908
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19705 5899 19763 5905
rect 19705 5896 19717 5899
rect 19300 5868 19717 5896
rect 19300 5856 19306 5868
rect 19705 5865 19717 5868
rect 19751 5865 19763 5899
rect 19705 5859 19763 5865
rect 23290 5856 23296 5908
rect 23348 5896 23354 5908
rect 23477 5899 23535 5905
rect 23477 5896 23489 5899
rect 23348 5868 23489 5896
rect 23348 5856 23354 5868
rect 23477 5865 23489 5868
rect 23523 5865 23535 5899
rect 23477 5859 23535 5865
rect 11149 5831 11207 5837
rect 11149 5828 11161 5831
rect 10704 5800 11161 5828
rect 4982 5720 4988 5772
rect 5040 5720 5046 5772
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5629 5695 5687 5701
rect 5629 5692 5641 5695
rect 5592 5664 5641 5692
rect 5592 5652 5598 5664
rect 5629 5661 5641 5664
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 10594 5652 10600 5704
rect 10652 5692 10658 5704
rect 10704 5701 10732 5800
rect 11149 5797 11161 5800
rect 11195 5797 11207 5831
rect 14274 5828 14280 5840
rect 11149 5791 11207 5797
rect 13188 5800 14280 5828
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 10870 5760 10876 5772
rect 10827 5732 10876 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10652 5664 10701 5692
rect 10652 5652 10658 5664
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10888 5692 10916 5720
rect 11333 5695 11391 5701
rect 11333 5692 11345 5695
rect 10888 5664 11345 5692
rect 10689 5655 10747 5661
rect 11333 5661 11345 5664
rect 11379 5661 11391 5695
rect 11333 5655 11391 5661
rect 12862 5695 12920 5701
rect 12862 5661 12874 5695
rect 12908 5692 12920 5695
rect 13188 5692 13216 5800
rect 14274 5788 14280 5800
rect 14332 5788 14338 5840
rect 18966 5788 18972 5840
rect 19024 5828 19030 5840
rect 19024 5800 19288 5828
rect 19024 5788 19030 5800
rect 13262 5720 13268 5772
rect 13320 5760 13326 5772
rect 13725 5763 13783 5769
rect 13725 5760 13737 5763
rect 13320 5732 13737 5760
rect 13320 5720 13326 5732
rect 13725 5729 13737 5732
rect 13771 5729 13783 5763
rect 13725 5723 13783 5729
rect 13909 5763 13967 5769
rect 13909 5729 13921 5763
rect 13955 5760 13967 5763
rect 14366 5760 14372 5772
rect 13955 5732 14372 5760
rect 13955 5729 13967 5732
rect 13909 5723 13967 5729
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 17681 5763 17739 5769
rect 17681 5729 17693 5763
rect 17727 5760 17739 5763
rect 18046 5760 18052 5772
rect 17727 5732 18052 5760
rect 17727 5729 17739 5732
rect 17681 5723 17739 5729
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 19260 5769 19288 5800
rect 19061 5763 19119 5769
rect 19061 5729 19073 5763
rect 19107 5729 19119 5763
rect 19061 5723 19119 5729
rect 19245 5763 19303 5769
rect 19245 5729 19257 5763
rect 19291 5729 19303 5763
rect 19613 5763 19671 5769
rect 19613 5760 19625 5763
rect 19245 5723 19303 5729
rect 19352 5732 19625 5760
rect 12908 5664 13216 5692
rect 12908 5661 12920 5664
rect 12862 5655 12920 5661
rect 13446 5652 13452 5704
rect 13504 5652 13510 5704
rect 17586 5652 17592 5704
rect 17644 5652 17650 5704
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 19076 5692 19104 5723
rect 19352 5692 19380 5732
rect 19613 5729 19625 5732
rect 19659 5760 19671 5763
rect 19659 5732 20024 5760
rect 19659 5729 19671 5732
rect 19613 5723 19671 5729
rect 19996 5704 20024 5732
rect 19076 5664 19380 5692
rect 19429 5695 19487 5701
rect 18877 5655 18935 5661
rect 19429 5661 19441 5695
rect 19475 5692 19487 5695
rect 19475 5664 19932 5692
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 13265 5627 13323 5633
rect 13265 5593 13277 5627
rect 13311 5624 13323 5627
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 13311 5596 13553 5624
rect 13311 5593 13323 5596
rect 13265 5587 13323 5593
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 18892 5624 18920 5655
rect 19444 5624 19472 5655
rect 19904 5633 19932 5664
rect 19978 5652 19984 5704
rect 20036 5692 20042 5704
rect 20073 5695 20131 5701
rect 20073 5692 20085 5695
rect 20036 5664 20085 5692
rect 20036 5652 20042 5664
rect 20073 5661 20085 5664
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 23382 5652 23388 5704
rect 23440 5692 23446 5704
rect 23661 5695 23719 5701
rect 23661 5692 23673 5695
rect 23440 5664 23673 5692
rect 23440 5652 23446 5664
rect 23661 5661 23673 5664
rect 23707 5661 23719 5695
rect 23661 5655 23719 5661
rect 18892 5596 19472 5624
rect 19889 5627 19947 5633
rect 13541 5587 13599 5593
rect 19889 5593 19901 5627
rect 19935 5624 19947 5627
rect 20162 5624 20168 5636
rect 19935 5596 20168 5624
rect 19935 5593 19947 5596
rect 19889 5587 19947 5593
rect 20162 5584 20168 5596
rect 20220 5584 20226 5636
rect 5074 5516 5080 5568
rect 5132 5516 5138 5568
rect 5166 5516 5172 5568
rect 5224 5516 5230 5568
rect 11514 5516 11520 5568
rect 11572 5516 11578 5568
rect 13081 5559 13139 5565
rect 13081 5525 13093 5559
rect 13127 5556 13139 5559
rect 13814 5556 13820 5568
rect 13127 5528 13820 5556
rect 13127 5525 13139 5528
rect 13081 5519 13139 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 1104 5466 24012 5488
rect 1104 5414 4473 5466
rect 4525 5414 4537 5466
rect 4589 5414 4601 5466
rect 4653 5414 4665 5466
rect 4717 5414 4729 5466
rect 4781 5414 10200 5466
rect 10252 5414 10264 5466
rect 10316 5414 10328 5466
rect 10380 5414 10392 5466
rect 10444 5414 10456 5466
rect 10508 5414 15927 5466
rect 15979 5414 15991 5466
rect 16043 5414 16055 5466
rect 16107 5414 16119 5466
rect 16171 5414 16183 5466
rect 16235 5414 21654 5466
rect 21706 5414 21718 5466
rect 21770 5414 21782 5466
rect 21834 5414 21846 5466
rect 21898 5414 21910 5466
rect 21962 5414 24012 5466
rect 1104 5392 24012 5414
rect 5074 5312 5080 5364
rect 5132 5312 5138 5364
rect 5534 5312 5540 5364
rect 5592 5312 5598 5364
rect 14366 5312 14372 5364
rect 14424 5312 14430 5364
rect 14918 5312 14924 5364
rect 14976 5352 14982 5364
rect 19889 5355 19947 5361
rect 14976 5324 18552 5352
rect 14976 5312 14982 5324
rect 4985 5287 5043 5293
rect 4985 5253 4997 5287
rect 5031 5284 5043 5287
rect 5350 5284 5356 5296
rect 5031 5256 5356 5284
rect 5031 5253 5043 5256
rect 4985 5247 5043 5253
rect 5350 5244 5356 5256
rect 5408 5244 5414 5296
rect 10505 5287 10563 5293
rect 8036 5256 8800 5284
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4396 5188 4629 5216
rect 4396 5176 4402 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4798 5176 4804 5228
rect 4856 5176 4862 5228
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 4890 5108 4896 5160
rect 4948 5148 4954 5160
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 4948 5120 5641 5148
rect 4948 5108 4954 5120
rect 5629 5117 5641 5120
rect 5675 5117 5687 5151
rect 5629 5111 5687 5117
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 8036 5157 8064 5256
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8021 5151 8079 5157
rect 8021 5148 8033 5151
rect 7708 5120 8033 5148
rect 7708 5108 7714 5120
rect 8021 5117 8033 5120
rect 8067 5117 8079 5151
rect 8021 5111 8079 5117
rect 8128 5080 8156 5179
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8772 5157 8800 5256
rect 10505 5253 10517 5287
rect 10551 5284 10563 5287
rect 11514 5284 11520 5296
rect 10551 5256 11520 5284
rect 10551 5253 10563 5256
rect 10505 5247 10563 5253
rect 11514 5244 11520 5256
rect 11572 5244 11578 5296
rect 17773 5287 17831 5293
rect 17773 5253 17785 5287
rect 17819 5284 17831 5287
rect 18049 5287 18107 5293
rect 18049 5284 18061 5287
rect 17819 5256 18061 5284
rect 17819 5253 17831 5256
rect 17773 5247 17831 5253
rect 18049 5253 18061 5256
rect 18095 5253 18107 5287
rect 18049 5247 18107 5253
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 11330 5216 11336 5228
rect 10735 5188 11336 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 14734 5176 14740 5228
rect 14792 5176 14798 5228
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 8352 5120 8493 5148
rect 8352 5108 8358 5120
rect 8481 5117 8493 5120
rect 8527 5117 8539 5151
rect 8481 5111 8539 5117
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 14826 5108 14832 5160
rect 14884 5148 14890 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 14884 5120 15301 5148
rect 14884 5108 14890 5120
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 8941 5083 8999 5089
rect 8941 5080 8953 5083
rect 8128 5052 8953 5080
rect 8941 5049 8953 5052
rect 8987 5080 8999 5083
rect 10321 5083 10379 5089
rect 10321 5080 10333 5083
rect 8987 5052 10333 5080
rect 8987 5049 8999 5052
rect 8941 5043 8999 5049
rect 10321 5049 10333 5052
rect 10367 5049 10379 5083
rect 15396 5080 15424 5179
rect 17862 5176 17868 5228
rect 17920 5176 17926 5228
rect 15746 5108 15752 5160
rect 15804 5108 15810 5160
rect 17405 5151 17463 5157
rect 17405 5117 17417 5151
rect 17451 5148 17463 5151
rect 17494 5148 17500 5160
rect 17451 5120 17500 5148
rect 17451 5117 17463 5120
rect 17405 5111 17463 5117
rect 17494 5108 17500 5120
rect 17552 5108 17558 5160
rect 17589 5151 17647 5157
rect 17589 5117 17601 5151
rect 17635 5148 17647 5151
rect 18046 5148 18052 5160
rect 17635 5120 18052 5148
rect 17635 5117 17647 5120
rect 17589 5111 17647 5117
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 18233 5083 18291 5089
rect 18233 5080 18245 5083
rect 15396 5052 18245 5080
rect 10321 5043 10379 5049
rect 15764 5024 15792 5052
rect 18233 5049 18245 5052
rect 18279 5049 18291 5083
rect 18524 5080 18552 5324
rect 19889 5321 19901 5355
rect 19935 5352 19947 5355
rect 19978 5352 19984 5364
rect 19935 5324 19984 5352
rect 19935 5321 19947 5324
rect 19889 5315 19947 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20162 5312 20168 5364
rect 20220 5352 20226 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 20220 5324 20729 5352
rect 20220 5312 20226 5324
rect 20717 5321 20729 5324
rect 20763 5321 20775 5355
rect 20717 5315 20775 5321
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5216 20315 5219
rect 20806 5216 20812 5228
rect 20303 5188 20812 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5216 21143 5219
rect 21358 5216 21364 5228
rect 21131 5188 21364 5216
rect 21131 5185 21143 5188
rect 21085 5179 21143 5185
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 23658 5176 23664 5228
rect 23716 5176 23722 5228
rect 20346 5108 20352 5160
rect 20404 5108 20410 5160
rect 20438 5108 20444 5160
rect 20496 5108 20502 5160
rect 20898 5108 20904 5160
rect 20956 5148 20962 5160
rect 21177 5151 21235 5157
rect 21177 5148 21189 5151
rect 20956 5120 21189 5148
rect 20956 5108 20962 5120
rect 21177 5117 21189 5120
rect 21223 5117 21235 5151
rect 21177 5111 21235 5117
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5148 21327 5151
rect 21450 5148 21456 5160
rect 21315 5120 21456 5148
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 21450 5108 21456 5120
rect 21508 5148 21514 5160
rect 23106 5148 23112 5160
rect 21508 5120 23112 5148
rect 21508 5108 21514 5120
rect 23106 5108 23112 5120
rect 23164 5108 23170 5160
rect 23477 5083 23535 5089
rect 23477 5080 23489 5083
rect 18524 5052 23489 5080
rect 18233 5043 18291 5049
rect 23477 5049 23489 5052
rect 23523 5049 23535 5083
rect 23477 5043 23535 5049
rect 8570 4972 8576 5024
rect 8628 4972 8634 5024
rect 15746 4972 15752 5024
rect 15804 4972 15810 5024
rect 1104 4922 24012 4944
rect 1104 4870 3813 4922
rect 3865 4870 3877 4922
rect 3929 4870 3941 4922
rect 3993 4870 4005 4922
rect 4057 4870 4069 4922
rect 4121 4870 9540 4922
rect 9592 4870 9604 4922
rect 9656 4870 9668 4922
rect 9720 4870 9732 4922
rect 9784 4870 9796 4922
rect 9848 4870 15267 4922
rect 15319 4870 15331 4922
rect 15383 4870 15395 4922
rect 15447 4870 15459 4922
rect 15511 4870 15523 4922
rect 15575 4870 20994 4922
rect 21046 4870 21058 4922
rect 21110 4870 21122 4922
rect 21174 4870 21186 4922
rect 21238 4870 21250 4922
rect 21302 4870 24012 4922
rect 1104 4848 24012 4870
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 5537 4811 5595 4817
rect 5537 4808 5549 4811
rect 5500 4780 5549 4808
rect 5500 4768 5506 4780
rect 5537 4777 5549 4780
rect 5583 4777 5595 4811
rect 5537 4771 5595 4777
rect 10870 4768 10876 4820
rect 10928 4768 10934 4820
rect 11330 4768 11336 4820
rect 11388 4768 11394 4820
rect 14550 4768 14556 4820
rect 14608 4808 14614 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 14608 4780 14933 4808
rect 14608 4768 14614 4780
rect 14921 4777 14933 4780
rect 14967 4777 14979 4811
rect 14921 4771 14979 4777
rect 20346 4768 20352 4820
rect 20404 4808 20410 4820
rect 20898 4817 20904 4820
rect 20487 4811 20545 4817
rect 20487 4808 20499 4811
rect 20404 4780 20499 4808
rect 20404 4768 20410 4780
rect 20487 4777 20499 4780
rect 20533 4777 20545 4811
rect 20487 4771 20545 4777
rect 20855 4811 20904 4817
rect 20855 4777 20867 4811
rect 20901 4777 20904 4811
rect 20855 4771 20904 4777
rect 20898 4768 20904 4771
rect 20956 4768 20962 4820
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 7929 4743 7987 4749
rect 7929 4740 7941 4743
rect 7340 4712 7941 4740
rect 7340 4700 7346 4712
rect 7929 4709 7941 4712
rect 7975 4709 7987 4743
rect 15289 4743 15347 4749
rect 7929 4703 7987 4709
rect 10612 4712 11192 4740
rect 4890 4632 4896 4684
rect 4948 4632 4954 4684
rect 5810 4632 5816 4684
rect 5868 4632 5874 4684
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 5920 4644 7849 4672
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5920 4613 5948 4644
rect 7837 4641 7849 4644
rect 7883 4641 7895 4675
rect 8570 4672 8576 4684
rect 7837 4635 7895 4641
rect 8036 4644 8576 4672
rect 5905 4607 5963 4613
rect 5905 4604 5917 4607
rect 5684 4576 5917 4604
rect 5684 4564 5690 4576
rect 5905 4573 5917 4576
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 8036 4604 8064 4644
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 10612 4681 10640 4712
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 7699 4576 8064 4604
rect 8113 4607 8171 4613
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 8113 4573 8125 4607
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 10980 4604 11008 4635
rect 11164 4616 11192 4712
rect 15289 4709 15301 4743
rect 15335 4740 15347 4743
rect 15746 4740 15752 4752
rect 15335 4712 15752 4740
rect 15335 4709 15347 4712
rect 15289 4703 15347 4709
rect 15746 4700 15752 4712
rect 15804 4700 15810 4752
rect 21542 4632 21548 4684
rect 21600 4672 21606 4684
rect 22465 4675 22523 4681
rect 22465 4672 22477 4675
rect 21600 4644 22477 4672
rect 21600 4632 21606 4644
rect 22465 4641 22477 4644
rect 22511 4641 22523 4675
rect 22465 4635 22523 4641
rect 10551 4576 11008 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 4154 4496 4160 4548
rect 4212 4536 4218 4548
rect 5077 4539 5135 4545
rect 5077 4536 5089 4539
rect 4212 4508 5089 4536
rect 4212 4496 4218 4508
rect 5077 4505 5089 4508
rect 5123 4505 5135 4539
rect 5077 4499 5135 4505
rect 7466 4496 7472 4548
rect 7524 4496 7530 4548
rect 7558 4496 7564 4548
rect 7616 4536 7622 4548
rect 8128 4536 8156 4567
rect 10612 4548 10640 4576
rect 11146 4564 11152 4616
rect 11204 4564 11210 4616
rect 14826 4564 14832 4616
rect 14884 4604 14890 4616
rect 15105 4607 15163 4613
rect 15105 4604 15117 4607
rect 14884 4576 15117 4604
rect 14884 4564 14890 4576
rect 15105 4573 15117 4576
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 20590 4607 20648 4613
rect 20590 4573 20602 4607
rect 20636 4604 20648 4607
rect 20784 4607 20842 4613
rect 20636 4573 20668 4604
rect 20590 4567 20668 4573
rect 20784 4573 20796 4607
rect 20830 4604 20842 4607
rect 21358 4604 21364 4616
rect 20830 4576 21364 4604
rect 20830 4573 20842 4576
rect 20784 4567 20842 4573
rect 7616 4508 8156 4536
rect 7616 4496 7622 4508
rect 10594 4496 10600 4548
rect 10652 4496 10658 4548
rect 20640 4536 20668 4567
rect 21358 4564 21364 4576
rect 21416 4604 21422 4616
rect 23474 4604 23480 4616
rect 21416 4576 23480 4604
rect 21416 4564 21422 4576
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 23658 4564 23664 4616
rect 23716 4564 23722 4616
rect 20898 4536 20904 4548
rect 20640 4508 20904 4536
rect 20898 4496 20904 4508
rect 20956 4496 20962 4548
rect 4982 4428 4988 4480
rect 5040 4428 5046 4480
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 5224 4440 5457 4468
rect 5224 4428 5230 4440
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5445 4431 5503 4437
rect 8110 4428 8116 4480
rect 8168 4468 8174 4480
rect 8297 4471 8355 4477
rect 8297 4468 8309 4471
rect 8168 4440 8309 4468
rect 8168 4428 8174 4440
rect 8297 4437 8309 4440
rect 8343 4437 8355 4471
rect 8297 4431 8355 4437
rect 1104 4378 24012 4400
rect 1104 4326 4473 4378
rect 4525 4326 4537 4378
rect 4589 4326 4601 4378
rect 4653 4326 4665 4378
rect 4717 4326 4729 4378
rect 4781 4326 10200 4378
rect 10252 4326 10264 4378
rect 10316 4326 10328 4378
rect 10380 4326 10392 4378
rect 10444 4326 10456 4378
rect 10508 4326 15927 4378
rect 15979 4326 15991 4378
rect 16043 4326 16055 4378
rect 16107 4326 16119 4378
rect 16171 4326 16183 4378
rect 16235 4326 21654 4378
rect 21706 4326 21718 4378
rect 21770 4326 21782 4378
rect 21834 4326 21846 4378
rect 21898 4326 21910 4378
rect 21962 4326 24012 4378
rect 1104 4304 24012 4326
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 4525 4267 4583 4273
rect 4525 4264 4537 4267
rect 4396 4236 4537 4264
rect 4396 4224 4402 4236
rect 4525 4233 4537 4236
rect 4571 4233 4583 4267
rect 4525 4227 4583 4233
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 5261 4267 5319 4273
rect 5261 4264 5273 4267
rect 4856 4236 5273 4264
rect 4856 4224 4862 4236
rect 5261 4233 5273 4236
rect 5307 4233 5319 4267
rect 5261 4227 5319 4233
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7466 4264 7472 4276
rect 7055 4236 7472 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 8110 4224 8116 4276
rect 8168 4224 8174 4276
rect 11146 4264 11152 4276
rect 10060 4236 11152 4264
rect 10060 4205 10088 4236
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 18138 4224 18144 4276
rect 18196 4224 18202 4276
rect 10045 4199 10103 4205
rect 10045 4165 10057 4199
rect 10091 4165 10103 4199
rect 10045 4159 10103 4165
rect 10229 4199 10287 4205
rect 10229 4165 10241 4199
rect 10275 4196 10287 4199
rect 10594 4196 10600 4208
rect 10275 4168 10600 4196
rect 10275 4165 10287 4168
rect 10229 4159 10287 4165
rect 10594 4156 10600 4168
rect 10652 4156 10658 4208
rect 18156 4196 18184 4224
rect 15028 4168 16160 4196
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 4154 4128 4160 4140
rect 3743 4100 4160 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 4890 4128 4896 4140
rect 4847 4100 4896 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5184 4100 5457 4128
rect 5184 4069 5212 4100
rect 5445 4097 5457 4100
rect 5491 4128 5503 4131
rect 5810 4128 5816 4140
rect 5491 4100 5816 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 7282 4128 7288 4140
rect 6656 4100 7288 4128
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 3927 4032 4353 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 4341 4029 4353 4032
rect 4387 4060 4399 4063
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4387 4032 4721 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 4709 4029 4721 4032
rect 4755 4060 4767 4063
rect 5169 4063 5227 4069
rect 4755 4032 4844 4060
rect 4755 4029 4767 4032
rect 4709 4023 4767 4029
rect 4816 4004 4844 4032
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5626 4020 5632 4072
rect 5684 4020 5690 4072
rect 6656 4069 6684 4100
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 10686 4088 10692 4140
rect 10744 4088 10750 4140
rect 14369 4131 14427 4137
rect 14369 4097 14381 4131
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 6871 4032 7389 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7377 4029 7389 4032
rect 7423 4060 7435 4063
rect 7558 4060 7564 4072
rect 7423 4032 7564 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 7650 4020 7656 4072
rect 7708 4020 7714 4072
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7984 4032 8033 4060
rect 7984 4020 7990 4032
rect 8021 4029 8033 4032
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 9907 4032 10793 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 10873 4063 10931 4069
rect 10873 4029 10885 4063
rect 10919 4029 10931 4063
rect 10873 4023 10931 4029
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 4111 3964 4169 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 4157 3961 4169 3964
rect 4203 3961 4215 3995
rect 4157 3955 4215 3961
rect 4172 3924 4200 3955
rect 4798 3952 4804 4004
rect 4856 3952 4862 4004
rect 4890 3924 4896 3936
rect 4172 3896 4896 3924
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 7852 3924 7880 4020
rect 8478 3952 8484 4004
rect 8536 3952 8542 4004
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 10321 3995 10379 4001
rect 10321 3992 10333 3995
rect 10100 3964 10333 3992
rect 10100 3952 10106 3964
rect 10321 3961 10333 3964
rect 10367 3961 10379 3995
rect 10888 3992 10916 4023
rect 10321 3955 10379 3961
rect 10796 3964 10916 3992
rect 10796 3924 10824 3964
rect 7852 3896 10824 3924
rect 14384 3924 14412 4091
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4060 14795 4063
rect 14826 4060 14832 4072
rect 14783 4032 14832 4060
rect 14783 4029 14795 4032
rect 14737 4023 14795 4029
rect 14476 3992 14504 4023
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 15028 4069 15056 4168
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4128 15255 4131
rect 16025 4131 16083 4137
rect 16025 4128 16037 4131
rect 15243 4100 16037 4128
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 16025 4097 16037 4100
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 15102 4020 15108 4072
rect 15160 4020 15166 4072
rect 15838 4060 15844 4072
rect 15212 4032 15844 4060
rect 15212 3992 15240 4032
rect 15838 4020 15844 4032
rect 15896 4020 15902 4072
rect 16132 4060 16160 4168
rect 17972 4168 18184 4196
rect 17586 4088 17592 4140
rect 17644 4088 17650 4140
rect 17972 4128 18000 4168
rect 17880 4100 18000 4128
rect 16132 4032 17632 4060
rect 14476 3964 15240 3992
rect 15562 3952 15568 4004
rect 15620 3952 15626 4004
rect 15657 3995 15715 4001
rect 15657 3961 15669 3995
rect 15703 3961 15715 3995
rect 15657 3955 15715 3961
rect 14826 3924 14832 3936
rect 14384 3896 14832 3924
rect 14826 3884 14832 3896
rect 14884 3924 14890 3936
rect 15672 3924 15700 3955
rect 16666 3952 16672 4004
rect 16724 3992 16730 4004
rect 17221 3995 17279 4001
rect 17221 3992 17233 3995
rect 16724 3964 17233 3992
rect 16724 3952 16730 3964
rect 17221 3961 17233 3964
rect 17267 3961 17279 3995
rect 17604 3992 17632 4032
rect 17678 4020 17684 4072
rect 17736 4020 17742 4072
rect 17880 4069 17908 4100
rect 18138 4088 18144 4140
rect 18196 4128 18202 4140
rect 18417 4131 18475 4137
rect 18417 4128 18429 4131
rect 18196 4100 18429 4128
rect 18196 4088 18202 4100
rect 18417 4097 18429 4100
rect 18463 4097 18475 4131
rect 18417 4091 18475 4097
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4029 17923 4063
rect 17865 4023 17923 4029
rect 17880 3992 17908 4023
rect 18046 4020 18052 4072
rect 18104 4020 18110 4072
rect 18322 4020 18328 4072
rect 18380 4020 18386 4072
rect 17604 3964 17908 3992
rect 17221 3955 17279 3961
rect 14884 3896 15700 3924
rect 14884 3884 14890 3896
rect 1104 3834 24012 3856
rect 1104 3782 3813 3834
rect 3865 3782 3877 3834
rect 3929 3782 3941 3834
rect 3993 3782 4005 3834
rect 4057 3782 4069 3834
rect 4121 3782 9540 3834
rect 9592 3782 9604 3834
rect 9656 3782 9668 3834
rect 9720 3782 9732 3834
rect 9784 3782 9796 3834
rect 9848 3782 15267 3834
rect 15319 3782 15331 3834
rect 15383 3782 15395 3834
rect 15447 3782 15459 3834
rect 15511 3782 15523 3834
rect 15575 3782 20994 3834
rect 21046 3782 21058 3834
rect 21110 3782 21122 3834
rect 21174 3782 21186 3834
rect 21238 3782 21250 3834
rect 21302 3782 24012 3834
rect 1104 3760 24012 3782
rect 4982 3680 4988 3732
rect 5040 3680 5046 3732
rect 7926 3680 7932 3732
rect 7984 3680 7990 3732
rect 10594 3680 10600 3732
rect 10652 3680 10658 3732
rect 10686 3680 10692 3732
rect 10744 3680 10750 3732
rect 14734 3680 14740 3732
rect 14792 3680 14798 3732
rect 15194 3680 15200 3732
rect 15252 3680 15258 3732
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 17586 3720 17592 3732
rect 16899 3692 17592 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 17678 3680 17684 3732
rect 17736 3720 17742 3732
rect 17773 3723 17831 3729
rect 17773 3720 17785 3723
rect 17736 3692 17785 3720
rect 17736 3680 17742 3692
rect 17773 3689 17785 3692
rect 17819 3689 17831 3723
rect 17773 3683 17831 3689
rect 18322 3680 18328 3732
rect 18380 3680 18386 3732
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 23477 3723 23535 3729
rect 23477 3720 23489 3723
rect 20956 3692 23489 3720
rect 20956 3680 20962 3692
rect 23477 3689 23489 3692
rect 23523 3689 23535 3723
rect 23477 3683 23535 3689
rect 10612 3652 10640 3680
rect 11057 3655 11115 3661
rect 11057 3652 11069 3655
rect 10612 3624 11069 3652
rect 11057 3621 11069 3624
rect 11103 3621 11115 3655
rect 11057 3615 11115 3621
rect 11517 3655 11575 3661
rect 11517 3621 11529 3655
rect 11563 3621 11575 3655
rect 12526 3652 12532 3664
rect 11517 3615 11575 3621
rect 11624 3624 12532 3652
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 11146 3584 11152 3596
rect 10919 3556 11152 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4890 3516 4896 3528
rect 4663 3488 4896 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7282 3516 7288 3528
rect 6972 3488 7288 3516
rect 6972 3476 6978 3488
rect 7282 3476 7288 3488
rect 7340 3516 7346 3528
rect 7561 3519 7619 3525
rect 7561 3516 7573 3519
rect 7340 3488 7573 3516
rect 7340 3476 7346 3488
rect 7561 3485 7573 3488
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7708 3488 7757 3516
rect 7708 3476 7714 3488
rect 7745 3485 7757 3488
rect 7791 3485 7803 3519
rect 10060 3516 10088 3547
rect 11146 3544 11152 3556
rect 11204 3584 11210 3596
rect 11532 3584 11560 3615
rect 11204 3556 11560 3584
rect 11204 3544 11210 3556
rect 11624 3516 11652 3624
rect 12526 3612 12532 3624
rect 12584 3652 12590 3664
rect 13722 3652 13728 3664
rect 12584 3624 13728 3652
rect 12584 3612 12590 3624
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 17221 3655 17279 3661
rect 17221 3621 17233 3655
rect 17267 3652 17279 3655
rect 17313 3655 17371 3661
rect 17313 3652 17325 3655
rect 17267 3624 17325 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17313 3621 17325 3624
rect 17359 3652 17371 3655
rect 18138 3652 18144 3664
rect 17359 3624 18144 3652
rect 17359 3621 17371 3624
rect 17313 3615 17371 3621
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 12066 3544 12072 3596
rect 12124 3544 12130 3596
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3584 14427 3587
rect 14826 3584 14832 3596
rect 14415 3556 14832 3584
rect 14415 3553 14427 3556
rect 14369 3547 14427 3553
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 17681 3587 17739 3593
rect 17681 3553 17693 3587
rect 17727 3584 17739 3587
rect 17862 3584 17868 3596
rect 17727 3556 17868 3584
rect 17727 3553 17739 3556
rect 17681 3547 17739 3553
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 12462 3519 12520 3525
rect 12462 3516 12474 3519
rect 10060 3488 11652 3516
rect 11900 3488 12474 3516
rect 7745 3479 7803 3485
rect 4798 3408 4804 3460
rect 4856 3408 4862 3460
rect 9858 3408 9864 3460
rect 9916 3448 9922 3460
rect 10229 3451 10287 3457
rect 10229 3448 10241 3451
rect 9916 3420 10241 3448
rect 9916 3408 9922 3420
rect 10229 3417 10241 3420
rect 10275 3417 10287 3451
rect 10229 3411 10287 3417
rect 11900 3392 11928 3488
rect 12462 3485 12474 3488
rect 12508 3485 12520 3519
rect 12462 3479 12520 3485
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3516 14611 3519
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14599 3488 15025 3516
rect 14599 3485 14611 3488
rect 14553 3479 14611 3485
rect 15013 3485 15025 3488
rect 15059 3516 15071 3519
rect 15838 3516 15844 3528
rect 15059 3488 15844 3516
rect 15059 3485 15071 3488
rect 15013 3479 15071 3485
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 17497 3519 17555 3525
rect 17497 3516 17509 3519
rect 17083 3488 17509 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 17497 3485 17509 3488
rect 17543 3516 17555 3519
rect 17957 3519 18015 3525
rect 17957 3516 17969 3519
rect 17543 3488 17969 3516
rect 17543 3485 17555 3488
rect 17497 3479 17555 3485
rect 17957 3485 17969 3488
rect 18003 3516 18015 3519
rect 18340 3516 18368 3680
rect 18969 3587 19027 3593
rect 18969 3553 18981 3587
rect 19015 3584 19027 3587
rect 21450 3584 21456 3596
rect 19015 3556 21456 3584
rect 19015 3553 19027 3556
rect 18969 3547 19027 3553
rect 18984 3516 19012 3547
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 18003 3488 18368 3516
rect 18432 3488 19012 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 14826 3408 14832 3460
rect 14884 3408 14890 3460
rect 18138 3408 18144 3460
rect 18196 3408 18202 3460
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 18432 3448 18460 3488
rect 23658 3476 23664 3528
rect 23716 3476 23722 3528
rect 18288 3420 18460 3448
rect 18693 3451 18751 3457
rect 18288 3408 18294 3420
rect 18693 3417 18705 3451
rect 18739 3448 18751 3451
rect 19518 3448 19524 3460
rect 18739 3420 19524 3448
rect 18739 3417 18751 3420
rect 18693 3411 18751 3417
rect 19518 3408 19524 3420
rect 19576 3408 19582 3460
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10137 3383 10195 3389
rect 10137 3380 10149 3383
rect 10100 3352 10149 3380
rect 10100 3340 10106 3352
rect 10137 3349 10149 3352
rect 10183 3349 10195 3383
rect 10137 3343 10195 3349
rect 11882 3340 11888 3392
rect 11940 3340 11946 3392
rect 11977 3383 12035 3389
rect 11977 3349 11989 3383
rect 12023 3380 12035 3383
rect 12391 3383 12449 3389
rect 12391 3380 12403 3383
rect 12023 3352 12403 3380
rect 12023 3349 12035 3352
rect 11977 3343 12035 3349
rect 12391 3349 12403 3352
rect 12437 3349 12449 3383
rect 12391 3343 12449 3349
rect 18782 3340 18788 3392
rect 18840 3340 18846 3392
rect 1104 3290 24012 3312
rect 1104 3238 4473 3290
rect 4525 3238 4537 3290
rect 4589 3238 4601 3290
rect 4653 3238 4665 3290
rect 4717 3238 4729 3290
rect 4781 3238 10200 3290
rect 10252 3238 10264 3290
rect 10316 3238 10328 3290
rect 10380 3238 10392 3290
rect 10444 3238 10456 3290
rect 10508 3238 15927 3290
rect 15979 3238 15991 3290
rect 16043 3238 16055 3290
rect 16107 3238 16119 3290
rect 16171 3238 16183 3290
rect 16235 3238 21654 3290
rect 21706 3238 21718 3290
rect 21770 3238 21782 3290
rect 21834 3238 21846 3290
rect 21898 3238 21910 3290
rect 21962 3238 24012 3290
rect 1104 3216 24012 3238
rect 4798 3136 4804 3188
rect 4856 3136 4862 3188
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 6914 3176 6920 3188
rect 6687 3148 6920 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7009 3179 7067 3185
rect 7009 3145 7021 3179
rect 7055 3176 7067 3179
rect 7374 3176 7380 3188
rect 7055 3148 7380 3176
rect 7055 3145 7067 3148
rect 7009 3139 7067 3145
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 7469 3179 7527 3185
rect 7469 3145 7481 3179
rect 7515 3176 7527 3179
rect 7650 3176 7656 3188
rect 7515 3148 7656 3176
rect 7515 3145 7527 3148
rect 7469 3139 7527 3145
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10275 3179 10333 3185
rect 10275 3176 10287 3179
rect 10100 3148 10287 3176
rect 10100 3136 10106 3148
rect 10275 3145 10287 3148
rect 10321 3145 10333 3179
rect 10275 3139 10333 3145
rect 14645 3179 14703 3185
rect 14645 3145 14657 3179
rect 14691 3176 14703 3179
rect 14826 3176 14832 3188
rect 14691 3148 14832 3176
rect 14691 3145 14703 3148
rect 14645 3139 14703 3145
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 15473 3179 15531 3185
rect 15473 3145 15485 3179
rect 15519 3176 15531 3179
rect 15838 3176 15844 3188
rect 15519 3148 15844 3176
rect 15519 3145 15531 3148
rect 15473 3139 15531 3145
rect 15838 3136 15844 3148
rect 15896 3136 15902 3188
rect 17681 3179 17739 3185
rect 15948 3148 16160 3176
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 5169 3111 5227 3117
rect 5169 3108 5181 3111
rect 4212 3080 5181 3108
rect 4212 3068 4218 3080
rect 5169 3077 5181 3080
rect 5215 3108 5227 3111
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 5215 3080 5856 3108
rect 5215 3077 5227 3080
rect 5169 3071 5227 3077
rect 4522 3000 4528 3052
rect 4580 3049 4586 3052
rect 5828 3049 5856 3080
rect 6932 3080 7849 3108
rect 6932 3052 6960 3080
rect 7837 3077 7849 3080
rect 7883 3108 7895 3111
rect 12066 3108 12072 3120
rect 7883 3080 8524 3108
rect 7883 3077 7895 3080
rect 7837 3071 7895 3077
rect 4580 3043 4618 3049
rect 4606 3009 4618 3043
rect 4580 3003 4618 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 5675 3043 5733 3049
rect 5675 3040 5687 3043
rect 5307 3012 5687 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 5675 3009 5687 3012
rect 5721 3009 5733 3043
rect 5675 3003 5733 3009
rect 5778 3043 5856 3049
rect 5778 3009 5790 3043
rect 5824 3012 5856 3043
rect 5824 3009 5836 3012
rect 5778 3003 5836 3009
rect 4580 3000 4586 3003
rect 6914 3000 6920 3052
rect 6972 3000 6978 3052
rect 8496 3049 8524 3080
rect 7929 3043 7987 3049
rect 7024 3012 7328 3040
rect 4246 2932 4252 2984
rect 4304 2972 4310 2984
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 4304 2944 5365 2972
rect 4304 2932 4310 2944
rect 5353 2941 5365 2944
rect 5399 2972 5411 2975
rect 7024 2972 7052 3012
rect 5399 2944 7052 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 7098 2932 7104 2984
rect 7156 2932 7162 2984
rect 7190 2932 7196 2984
rect 7248 2932 7254 2984
rect 7300 2972 7328 3012
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 8343 3043 8401 3049
rect 8343 3040 8355 3043
rect 7975 3012 8355 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8343 3009 8355 3012
rect 8389 3009 8401 3043
rect 8343 3003 8401 3009
rect 8446 3043 8524 3049
rect 8446 3009 8458 3043
rect 8492 3012 8524 3043
rect 9048 3080 12072 3108
rect 8492 3009 8504 3012
rect 8446 3003 8504 3009
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7300 2944 8033 2972
rect 8021 2941 8033 2944
rect 8067 2972 8079 2975
rect 9048 2972 9076 3080
rect 12066 3068 12072 3080
rect 12124 3108 12130 3120
rect 15948 3108 15976 3148
rect 12124 3080 15976 3108
rect 12124 3068 12130 3080
rect 14660 3052 14688 3080
rect 16022 3068 16028 3120
rect 16080 3068 16086 3120
rect 9858 3040 9864 3052
rect 8067 2944 9076 2972
rect 9140 3012 9864 3040
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 9140 2904 9168 3012
rect 9858 3000 9864 3012
rect 9916 3040 9922 3052
rect 10172 3043 10230 3049
rect 10172 3040 10184 3043
rect 9916 3012 10184 3040
rect 9916 3000 9922 3012
rect 10172 3009 10184 3012
rect 10218 3009 10230 3043
rect 10172 3003 10230 3009
rect 14642 3000 14648 3052
rect 14700 3000 14706 3052
rect 15010 3000 15016 3052
rect 15068 3000 15074 3052
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 15841 3043 15899 3049
rect 15841 3040 15853 3043
rect 15712 3012 15853 3040
rect 15712 3000 15718 3012
rect 15841 3009 15853 3012
rect 15887 3040 15899 3043
rect 16040 3040 16068 3068
rect 15887 3012 16068 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 15102 2932 15108 2984
rect 15160 2932 15166 2984
rect 15289 2975 15347 2981
rect 15289 2941 15301 2975
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 6886 2876 9168 2904
rect 6886 2848 6914 2876
rect 13722 2864 13728 2916
rect 13780 2904 13786 2916
rect 15304 2904 15332 2935
rect 15930 2932 15936 2984
rect 15988 2932 15994 2984
rect 16132 2981 16160 3148
rect 17681 3145 17693 3179
rect 17727 3176 17739 3179
rect 18138 3176 18144 3188
rect 17727 3148 18144 3176
rect 17727 3145 17739 3148
rect 17681 3139 17739 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 18782 3136 18788 3188
rect 18840 3185 18846 3188
rect 18840 3179 18889 3185
rect 18840 3145 18843 3179
rect 18877 3145 18889 3179
rect 18840 3139 18889 3145
rect 18840 3136 18846 3139
rect 23474 3136 23480 3188
rect 23532 3136 23538 3188
rect 18049 3111 18107 3117
rect 18049 3077 18061 3111
rect 18095 3108 18107 3111
rect 18095 3080 18736 3108
rect 18095 3077 18107 3080
rect 18049 3071 18107 3077
rect 18708 3049 18736 3080
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3040 18199 3043
rect 18555 3043 18613 3049
rect 18555 3040 18567 3043
rect 18187 3012 18567 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 18555 3009 18567 3012
rect 18601 3009 18613 3043
rect 18555 3003 18613 3009
rect 18658 3043 18736 3049
rect 18658 3009 18670 3043
rect 18704 3009 18736 3043
rect 18658 3003 18736 3009
rect 18934 3043 18992 3049
rect 18934 3009 18946 3043
rect 18980 3040 18992 3043
rect 19518 3040 19524 3052
rect 18980 3012 19524 3040
rect 18980 3009 18992 3012
rect 18934 3003 18992 3009
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2972 16175 2975
rect 18230 2972 18236 2984
rect 16163 2944 18236 2972
rect 16163 2941 16175 2944
rect 16117 2935 16175 2941
rect 18230 2932 18236 2944
rect 18288 2932 18294 2984
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2941 18383 2975
rect 18708 2972 18736 3003
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 23658 3000 23664 3052
rect 23716 3000 23722 3052
rect 19426 2972 19432 2984
rect 18708 2944 19432 2972
rect 18325 2935 18383 2941
rect 18340 2904 18368 2935
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 20438 2904 20444 2916
rect 13780 2876 20444 2904
rect 13780 2864 13786 2876
rect 20438 2864 20444 2876
rect 20496 2864 20502 2916
rect 4706 2845 4712 2848
rect 4663 2839 4712 2845
rect 4663 2805 4675 2839
rect 4709 2805 4712 2839
rect 4663 2799 4712 2805
rect 4706 2796 4712 2799
rect 4764 2796 4770 2848
rect 6822 2796 6828 2848
rect 6880 2808 6914 2848
rect 6880 2796 6886 2808
rect 15010 2796 15016 2848
rect 15068 2836 15074 2848
rect 17494 2836 17500 2848
rect 15068 2808 17500 2836
rect 15068 2796 15074 2808
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 1104 2746 24012 2768
rect 1104 2694 3813 2746
rect 3865 2694 3877 2746
rect 3929 2694 3941 2746
rect 3993 2694 4005 2746
rect 4057 2694 4069 2746
rect 4121 2694 9540 2746
rect 9592 2694 9604 2746
rect 9656 2694 9668 2746
rect 9720 2694 9732 2746
rect 9784 2694 9796 2746
rect 9848 2694 15267 2746
rect 15319 2694 15331 2746
rect 15383 2694 15395 2746
rect 15447 2694 15459 2746
rect 15511 2694 15523 2746
rect 15575 2694 20994 2746
rect 21046 2694 21058 2746
rect 21110 2694 21122 2746
rect 21174 2694 21186 2746
rect 21238 2694 21250 2746
rect 21302 2694 24012 2746
rect 1104 2672 24012 2694
rect 4154 2592 4160 2644
rect 4212 2592 4218 2644
rect 4522 2592 4528 2644
rect 4580 2592 4586 2644
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 4890 2632 4896 2644
rect 4663 2604 4896 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6914 2632 6920 2644
rect 6135 2604 6920 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7423 2635 7481 2641
rect 7423 2632 7435 2635
rect 7156 2604 7435 2632
rect 7156 2592 7162 2604
rect 7423 2601 7435 2604
rect 7469 2601 7481 2635
rect 7423 2595 7481 2601
rect 10597 2635 10655 2641
rect 10597 2601 10609 2635
rect 10643 2632 10655 2635
rect 10962 2632 10968 2644
rect 10643 2604 10968 2632
rect 10643 2601 10655 2604
rect 10597 2595 10655 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 11882 2592 11888 2644
rect 11940 2592 11946 2644
rect 12529 2635 12587 2641
rect 12529 2601 12541 2635
rect 12575 2632 12587 2635
rect 12618 2632 12624 2644
rect 12575 2604 12624 2632
rect 12575 2601 12587 2604
rect 12529 2595 12587 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 13354 2632 13360 2644
rect 13219 2604 13360 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 14274 2592 14280 2644
rect 14332 2592 14338 2644
rect 14967 2635 15025 2641
rect 14967 2601 14979 2635
rect 15013 2632 15025 2635
rect 15102 2632 15108 2644
rect 15013 2604 15108 2632
rect 15013 2601 15025 2604
rect 14967 2595 15025 2601
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 15335 2635 15393 2641
rect 15335 2601 15347 2635
rect 15381 2632 15393 2635
rect 15930 2632 15936 2644
rect 15381 2604 15936 2632
rect 15381 2601 15393 2604
rect 15335 2595 15393 2601
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16022 2592 16028 2644
rect 16080 2632 16086 2644
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 16080 2604 18797 2632
rect 16080 2592 16086 2604
rect 18785 2601 18797 2604
rect 18831 2601 18843 2635
rect 18785 2595 18843 2601
rect 19426 2592 19432 2644
rect 19484 2592 19490 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 19576 2604 21373 2632
rect 19576 2592 19582 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 6822 2564 6828 2576
rect 5675 2536 6828 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 6822 2524 6828 2536
rect 6880 2524 6886 2576
rect 7282 2524 7288 2576
rect 7340 2524 7346 2576
rect 15473 2567 15531 2573
rect 15473 2533 15485 2567
rect 15519 2564 15531 2567
rect 16482 2564 16488 2576
rect 15519 2536 16488 2564
rect 15519 2533 15531 2536
rect 15473 2527 15531 2533
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 17494 2524 17500 2576
rect 17552 2524 17558 2576
rect 4706 2456 4712 2508
rect 4764 2496 4770 2508
rect 5077 2499 5135 2505
rect 5077 2496 5089 2499
rect 4764 2468 5089 2496
rect 4764 2456 4770 2468
rect 5077 2465 5089 2468
rect 5123 2465 5135 2499
rect 5077 2459 5135 2465
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 7190 2496 7196 2508
rect 5316 2468 7196 2496
rect 5316 2456 5322 2468
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3292 2400 3341 2428
rect 3292 2388 3298 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4338 2388 4344 2440
rect 4396 2388 4402 2440
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 4580 2400 4997 2428
rect 4580 2388 4586 2400
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 4985 2391 5043 2397
rect 5184 2400 5457 2428
rect 5184 2372 5212 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5868 2400 5917 2428
rect 5868 2388 5874 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7006 2428 7012 2440
rect 6779 2400 7012 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 7300 2428 7328 2524
rect 7494 2431 7552 2437
rect 7494 2428 7506 2431
rect 7300 2400 7506 2428
rect 7494 2397 7506 2400
rect 7540 2397 7552 2431
rect 7494 2391 7552 2397
rect 8018 2388 8024 2440
rect 8076 2388 8082 2440
rect 8662 2388 8668 2440
rect 8720 2388 8726 2440
rect 9306 2388 9312 2440
rect 9364 2388 9370 2440
rect 9950 2388 9956 2440
rect 10008 2388 10014 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10594 2428 10600 2440
rect 10459 2400 10600 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 11020 2400 11069 2428
rect 11020 2388 11026 2400
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12952 2400 13001 2428
rect 12952 2388 12958 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 14240 2400 14473 2428
rect 14240 2388 14246 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 15010 2388 15016 2440
rect 15068 2437 15074 2440
rect 15068 2431 15096 2437
rect 15084 2397 15096 2431
rect 15068 2391 15096 2397
rect 15264 2431 15322 2437
rect 15264 2397 15276 2431
rect 15310 2428 15322 2431
rect 15562 2428 15568 2440
rect 15310 2400 15568 2428
rect 15310 2397 15322 2400
rect 15264 2391 15322 2397
rect 15068 2388 15074 2391
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 5166 2320 5172 2372
rect 5224 2320 5230 2372
rect 10778 2360 10784 2372
rect 5276 2332 10784 2360
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 5276 2292 5304 2332
rect 10778 2320 10784 2332
rect 10836 2320 10842 2372
rect 14826 2320 14832 2372
rect 14884 2360 14890 2372
rect 15672 2360 15700 2391
rect 15838 2388 15844 2440
rect 15896 2428 15902 2440
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 15896 2400 15945 2428
rect 15896 2388 15902 2400
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16390 2388 16396 2440
rect 16448 2388 16454 2440
rect 17034 2388 17040 2440
rect 17092 2388 17098 2440
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17460 2400 17693 2428
rect 17460 2388 17466 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18012 2400 18337 2428
rect 18012 2388 18018 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 18969 2431 19027 2437
rect 18969 2428 18981 2431
rect 18748 2400 18981 2428
rect 18748 2388 18754 2400
rect 18969 2397 18981 2400
rect 19015 2397 19027 2431
rect 18969 2391 19027 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20254 2388 20260 2440
rect 20312 2388 20318 2440
rect 20806 2388 20812 2440
rect 20864 2428 20870 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20864 2400 20913 2428
rect 20864 2388 20870 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 21545 2431 21603 2437
rect 21545 2428 21557 2431
rect 21324 2400 21557 2428
rect 21324 2388 21330 2400
rect 21545 2397 21557 2400
rect 21591 2397 21603 2431
rect 21545 2391 21603 2397
rect 14884 2332 15700 2360
rect 14884 2320 14890 2332
rect 3559 2264 5304 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6512 2264 6561 2292
rect 6512 2252 6518 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 7837 2295 7895 2301
rect 7837 2292 7849 2295
rect 7800 2264 7849 2292
rect 7800 2252 7806 2264
rect 7837 2261 7849 2264
rect 7883 2261 7895 2295
rect 7837 2255 7895 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8444 2264 8493 2292
rect 8444 2252 8450 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 9088 2264 9137 2292
rect 9088 2252 9094 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9732 2264 9781 2292
rect 9732 2252 9738 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13596 2264 13645 2292
rect 13596 2252 13602 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15620 2264 15761 2292
rect 15620 2252 15626 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 16209 2295 16267 2301
rect 16209 2261 16221 2295
rect 16255 2292 16267 2295
rect 16298 2292 16304 2304
rect 16255 2264 16304 2292
rect 16255 2261 16267 2264
rect 16209 2255 16267 2261
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16816 2264 16865 2292
rect 16816 2252 16822 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18141 2295 18199 2301
rect 18141 2292 18153 2295
rect 18104 2264 18153 2292
rect 18104 2252 18110 2264
rect 18141 2261 18153 2264
rect 18187 2261 18199 2295
rect 18141 2255 18199 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 20036 2264 20085 2292
rect 20036 2252 20042 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20717 2295 20775 2301
rect 20717 2292 20729 2295
rect 20680 2264 20729 2292
rect 20680 2252 20686 2264
rect 20717 2261 20729 2264
rect 20763 2261 20775 2295
rect 20717 2255 20775 2261
rect 1104 2202 24012 2224
rect 1104 2150 4473 2202
rect 4525 2150 4537 2202
rect 4589 2150 4601 2202
rect 4653 2150 4665 2202
rect 4717 2150 4729 2202
rect 4781 2150 10200 2202
rect 10252 2150 10264 2202
rect 10316 2150 10328 2202
rect 10380 2150 10392 2202
rect 10444 2150 10456 2202
rect 10508 2150 15927 2202
rect 15979 2150 15991 2202
rect 16043 2150 16055 2202
rect 16107 2150 16119 2202
rect 16171 2150 16183 2202
rect 16235 2150 21654 2202
rect 21706 2150 21718 2202
rect 21770 2150 21782 2202
rect 21834 2150 21846 2202
rect 21898 2150 21910 2202
rect 21962 2150 24012 2202
rect 1104 2128 24012 2150
<< via1 >>
rect 4473 24998 4525 25050
rect 4537 24998 4589 25050
rect 4601 24998 4653 25050
rect 4665 24998 4717 25050
rect 4729 24998 4781 25050
rect 10200 24998 10252 25050
rect 10264 24998 10316 25050
rect 10328 24998 10380 25050
rect 10392 24998 10444 25050
rect 10456 24998 10508 25050
rect 15927 24998 15979 25050
rect 15991 24998 16043 25050
rect 16055 24998 16107 25050
rect 16119 24998 16171 25050
rect 16183 24998 16235 25050
rect 21654 24998 21706 25050
rect 21718 24998 21770 25050
rect 21782 24998 21834 25050
rect 21846 24998 21898 25050
rect 21910 24998 21962 25050
rect 5816 24760 5868 24812
rect 6460 24760 6512 24812
rect 7104 24760 7156 24812
rect 7748 24760 7800 24812
rect 8668 24803 8720 24812
rect 8668 24769 8677 24803
rect 8677 24769 8711 24803
rect 8711 24769 8720 24803
rect 8668 24760 8720 24769
rect 9128 24760 9180 24812
rect 9864 24760 9916 24812
rect 10048 24760 10100 24812
rect 11060 24760 11112 24812
rect 11612 24760 11664 24812
rect 12256 24760 12308 24812
rect 12900 24760 12952 24812
rect 13544 24760 13596 24812
rect 14464 24803 14516 24812
rect 14464 24769 14473 24803
rect 14473 24769 14507 24803
rect 14507 24769 14516 24803
rect 14464 24760 14516 24769
rect 14832 24760 14884 24812
rect 15752 24803 15804 24812
rect 15752 24769 15761 24803
rect 15761 24769 15795 24803
rect 15795 24769 15804 24803
rect 15752 24760 15804 24769
rect 16396 24803 16448 24812
rect 16396 24769 16405 24803
rect 16405 24769 16439 24803
rect 16439 24769 16448 24803
rect 16396 24760 16448 24769
rect 16764 24760 16816 24812
rect 17408 24760 17460 24812
rect 18052 24760 18104 24812
rect 20628 24760 20680 24812
rect 23664 24803 23716 24812
rect 23664 24769 23673 24803
rect 23673 24769 23707 24803
rect 23707 24769 23716 24803
rect 23664 24760 23716 24769
rect 22744 24735 22796 24744
rect 22744 24701 22753 24735
rect 22753 24701 22787 24735
rect 22787 24701 22796 24735
rect 22744 24692 22796 24701
rect 8392 24624 8444 24676
rect 9036 24624 9088 24676
rect 9680 24624 9732 24676
rect 10600 24624 10652 24676
rect 10968 24624 11020 24676
rect 14188 24624 14240 24676
rect 15476 24624 15528 24676
rect 16304 24624 16356 24676
rect 6092 24599 6144 24608
rect 6092 24565 6101 24599
rect 6101 24565 6135 24599
rect 6135 24565 6144 24599
rect 6092 24556 6144 24565
rect 6736 24599 6788 24608
rect 6736 24565 6745 24599
rect 6745 24565 6779 24599
rect 6779 24565 6788 24599
rect 6736 24556 6788 24565
rect 7380 24599 7432 24608
rect 7380 24565 7389 24599
rect 7389 24565 7423 24599
rect 7423 24565 7432 24599
rect 7380 24556 7432 24565
rect 9312 24556 9364 24608
rect 11888 24599 11940 24608
rect 11888 24565 11897 24599
rect 11897 24565 11931 24599
rect 11931 24565 11940 24599
rect 11888 24556 11940 24565
rect 12532 24599 12584 24608
rect 12532 24565 12541 24599
rect 12541 24565 12575 24599
rect 12575 24565 12584 24599
rect 12532 24556 12584 24565
rect 12808 24556 12860 24608
rect 13636 24599 13688 24608
rect 13636 24565 13645 24599
rect 13645 24565 13679 24599
rect 13679 24565 13688 24599
rect 13636 24556 13688 24565
rect 14924 24599 14976 24608
rect 14924 24565 14933 24599
rect 14933 24565 14967 24599
rect 14967 24565 14976 24599
rect 14924 24556 14976 24565
rect 16856 24599 16908 24608
rect 16856 24565 16865 24599
rect 16865 24565 16899 24599
rect 16899 24565 16908 24599
rect 16856 24556 16908 24565
rect 17592 24556 17644 24608
rect 18328 24599 18380 24608
rect 18328 24565 18337 24599
rect 18337 24565 18371 24599
rect 18371 24565 18380 24599
rect 18328 24556 18380 24565
rect 20904 24599 20956 24608
rect 20904 24565 20913 24599
rect 20913 24565 20947 24599
rect 20947 24565 20956 24599
rect 20904 24556 20956 24565
rect 3813 24454 3865 24506
rect 3877 24454 3929 24506
rect 3941 24454 3993 24506
rect 4005 24454 4057 24506
rect 4069 24454 4121 24506
rect 9540 24454 9592 24506
rect 9604 24454 9656 24506
rect 9668 24454 9720 24506
rect 9732 24454 9784 24506
rect 9796 24454 9848 24506
rect 15267 24454 15319 24506
rect 15331 24454 15383 24506
rect 15395 24454 15447 24506
rect 15459 24454 15511 24506
rect 15523 24454 15575 24506
rect 20994 24454 21046 24506
rect 21058 24454 21110 24506
rect 21122 24454 21174 24506
rect 21186 24454 21238 24506
rect 21250 24454 21302 24506
rect 23020 24259 23072 24268
rect 23020 24225 23029 24259
rect 23029 24225 23063 24259
rect 23063 24225 23072 24259
rect 23020 24216 23072 24225
rect 7380 24148 7432 24200
rect 16856 24148 16908 24200
rect 23664 24191 23716 24200
rect 23664 24157 23673 24191
rect 23673 24157 23707 24191
rect 23707 24157 23716 24191
rect 23664 24148 23716 24157
rect 8392 24012 8444 24064
rect 15568 24012 15620 24064
rect 4473 23910 4525 23962
rect 4537 23910 4589 23962
rect 4601 23910 4653 23962
rect 4665 23910 4717 23962
rect 4729 23910 4781 23962
rect 10200 23910 10252 23962
rect 10264 23910 10316 23962
rect 10328 23910 10380 23962
rect 10392 23910 10444 23962
rect 10456 23910 10508 23962
rect 15927 23910 15979 23962
rect 15991 23910 16043 23962
rect 16055 23910 16107 23962
rect 16119 23910 16171 23962
rect 16183 23910 16235 23962
rect 21654 23910 21706 23962
rect 21718 23910 21770 23962
rect 21782 23910 21834 23962
rect 21846 23910 21898 23962
rect 21910 23910 21962 23962
rect 8392 23851 8444 23860
rect 8392 23817 8401 23851
rect 8401 23817 8435 23851
rect 8435 23817 8444 23851
rect 8392 23808 8444 23817
rect 9312 23851 9364 23860
rect 9312 23817 9321 23851
rect 9321 23817 9355 23851
rect 9355 23817 9364 23851
rect 9312 23808 9364 23817
rect 14924 23808 14976 23860
rect 15568 23851 15620 23860
rect 15568 23817 15577 23851
rect 15577 23817 15611 23851
rect 15611 23817 15620 23851
rect 15568 23808 15620 23817
rect 17592 23851 17644 23860
rect 17592 23817 17601 23851
rect 17601 23817 17635 23851
rect 17635 23817 17644 23851
rect 17592 23808 17644 23817
rect 7380 23740 7432 23792
rect 16856 23740 16908 23792
rect 12348 23672 12400 23724
rect 8300 23647 8352 23656
rect 8300 23613 8309 23647
rect 8309 23613 8343 23647
rect 8343 23613 8352 23647
rect 8300 23604 8352 23613
rect 8760 23604 8812 23656
rect 14740 23647 14792 23656
rect 14740 23613 14749 23647
rect 14749 23613 14783 23647
rect 14783 23613 14792 23647
rect 14740 23604 14792 23613
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 18328 23672 18380 23724
rect 23388 23672 23440 23724
rect 20628 23604 20680 23656
rect 12348 23536 12400 23588
rect 8852 23511 8904 23520
rect 8852 23477 8861 23511
rect 8861 23477 8895 23511
rect 8895 23477 8904 23511
rect 8852 23468 8904 23477
rect 9036 23468 9088 23520
rect 14280 23511 14332 23520
rect 14280 23477 14289 23511
rect 14289 23477 14323 23511
rect 14323 23477 14332 23511
rect 14280 23468 14332 23477
rect 15016 23468 15068 23520
rect 17040 23468 17092 23520
rect 18052 23468 18104 23520
rect 23848 23468 23900 23520
rect 3813 23366 3865 23418
rect 3877 23366 3929 23418
rect 3941 23366 3993 23418
rect 4005 23366 4057 23418
rect 4069 23366 4121 23418
rect 9540 23366 9592 23418
rect 9604 23366 9656 23418
rect 9668 23366 9720 23418
rect 9732 23366 9784 23418
rect 9796 23366 9848 23418
rect 15267 23366 15319 23418
rect 15331 23366 15383 23418
rect 15395 23366 15447 23418
rect 15459 23366 15511 23418
rect 15523 23366 15575 23418
rect 20994 23366 21046 23418
rect 21058 23366 21110 23418
rect 21122 23366 21174 23418
rect 21186 23366 21238 23418
rect 21250 23366 21302 23418
rect 14740 23264 14792 23316
rect 6828 23128 6880 23180
rect 15660 23128 15712 23180
rect 22744 23128 22796 23180
rect 6092 23060 6144 23112
rect 8852 23060 8904 23112
rect 9036 23060 9088 23112
rect 14924 23060 14976 23112
rect 18052 23060 18104 23112
rect 18328 22992 18380 23044
rect 6368 22967 6420 22976
rect 6368 22933 6377 22967
rect 6377 22933 6411 22967
rect 6411 22933 6420 22967
rect 6368 22924 6420 22933
rect 9496 22924 9548 22976
rect 17408 22967 17460 22976
rect 17408 22933 17417 22967
rect 17417 22933 17451 22967
rect 17451 22933 17460 22967
rect 17408 22924 17460 22933
rect 4473 22822 4525 22874
rect 4537 22822 4589 22874
rect 4601 22822 4653 22874
rect 4665 22822 4717 22874
rect 4729 22822 4781 22874
rect 10200 22822 10252 22874
rect 10264 22822 10316 22874
rect 10328 22822 10380 22874
rect 10392 22822 10444 22874
rect 10456 22822 10508 22874
rect 15927 22822 15979 22874
rect 15991 22822 16043 22874
rect 16055 22822 16107 22874
rect 16119 22822 16171 22874
rect 16183 22822 16235 22874
rect 21654 22822 21706 22874
rect 21718 22822 21770 22874
rect 21782 22822 21834 22874
rect 21846 22822 21898 22874
rect 21910 22822 21962 22874
rect 9496 22763 9548 22772
rect 9496 22729 9505 22763
rect 9505 22729 9539 22763
rect 9539 22729 9548 22763
rect 9496 22720 9548 22729
rect 11888 22720 11940 22772
rect 20904 22720 20956 22772
rect 6736 22584 6788 22636
rect 8852 22584 8904 22636
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 15016 22652 15068 22704
rect 5540 22516 5592 22568
rect 8300 22516 8352 22568
rect 9036 22516 9088 22568
rect 9220 22516 9272 22568
rect 9588 22559 9640 22568
rect 9588 22525 9597 22559
rect 9597 22525 9631 22559
rect 9631 22525 9640 22559
rect 9588 22516 9640 22525
rect 12348 22559 12400 22568
rect 12348 22525 12357 22559
rect 12357 22525 12391 22559
rect 12391 22525 12400 22559
rect 12348 22516 12400 22525
rect 14280 22559 14332 22568
rect 14280 22525 14289 22559
rect 14289 22525 14323 22559
rect 14323 22525 14332 22559
rect 14280 22516 14332 22525
rect 14924 22516 14976 22568
rect 17408 22584 17460 22636
rect 23664 22627 23716 22636
rect 23664 22593 23673 22627
rect 23673 22593 23707 22627
rect 23707 22593 23716 22627
rect 23664 22584 23716 22593
rect 16764 22516 16816 22568
rect 17040 22559 17092 22568
rect 17040 22525 17049 22559
rect 17049 22525 17083 22559
rect 17083 22525 17092 22559
rect 17040 22516 17092 22525
rect 20628 22559 20680 22568
rect 20628 22525 20637 22559
rect 20637 22525 20671 22559
rect 20671 22525 20680 22559
rect 20628 22516 20680 22525
rect 23020 22516 23072 22568
rect 8852 22448 8904 22500
rect 16672 22448 16724 22500
rect 17500 22448 17552 22500
rect 6460 22423 6512 22432
rect 6460 22389 6469 22423
rect 6469 22389 6503 22423
rect 6503 22389 6512 22423
rect 6460 22380 6512 22389
rect 8944 22423 8996 22432
rect 8944 22389 8953 22423
rect 8953 22389 8987 22423
rect 8987 22389 8996 22423
rect 8944 22380 8996 22389
rect 9036 22423 9088 22432
rect 9036 22389 9045 22423
rect 9045 22389 9079 22423
rect 9079 22389 9088 22423
rect 9036 22380 9088 22389
rect 9312 22380 9364 22432
rect 9588 22380 9640 22432
rect 9956 22380 10008 22432
rect 11980 22380 12032 22432
rect 14648 22423 14700 22432
rect 14648 22389 14657 22423
rect 14657 22389 14691 22423
rect 14691 22389 14700 22423
rect 14648 22380 14700 22389
rect 14740 22423 14792 22432
rect 14740 22389 14749 22423
rect 14749 22389 14783 22423
rect 14783 22389 14792 22423
rect 14740 22380 14792 22389
rect 17224 22380 17276 22432
rect 20904 22380 20956 22432
rect 23112 22380 23164 22432
rect 3813 22278 3865 22330
rect 3877 22278 3929 22330
rect 3941 22278 3993 22330
rect 4005 22278 4057 22330
rect 4069 22278 4121 22330
rect 9540 22278 9592 22330
rect 9604 22278 9656 22330
rect 9668 22278 9720 22330
rect 9732 22278 9784 22330
rect 9796 22278 9848 22330
rect 15267 22278 15319 22330
rect 15331 22278 15383 22330
rect 15395 22278 15447 22330
rect 15459 22278 15511 22330
rect 15523 22278 15575 22330
rect 20994 22278 21046 22330
rect 21058 22278 21110 22330
rect 21122 22278 21174 22330
rect 21186 22278 21238 22330
rect 21250 22278 21302 22330
rect 5908 22176 5960 22228
rect 6828 22176 6880 22228
rect 8760 22176 8812 22228
rect 8852 22108 8904 22160
rect 9404 22176 9456 22228
rect 15660 22176 15712 22228
rect 17408 22176 17460 22228
rect 9220 22040 9272 22092
rect 15016 22083 15068 22092
rect 15016 22049 15025 22083
rect 15025 22049 15059 22083
rect 15059 22049 15068 22083
rect 15016 22040 15068 22049
rect 15108 22040 15160 22092
rect 16580 22108 16632 22160
rect 16672 22040 16724 22092
rect 17500 22083 17552 22092
rect 17500 22049 17509 22083
rect 17509 22049 17543 22083
rect 17543 22049 17552 22083
rect 17500 22040 17552 22049
rect 17592 22040 17644 22092
rect 6368 21972 6420 22024
rect 12532 21972 12584 22024
rect 14648 21972 14700 22024
rect 14924 21972 14976 22024
rect 16580 22015 16632 22024
rect 16580 21981 16589 22015
rect 16589 21981 16623 22015
rect 16623 21981 16632 22015
rect 16580 21972 16632 21981
rect 6460 21947 6512 21956
rect 6460 21913 6469 21947
rect 6469 21913 6503 21947
rect 6503 21913 6512 21947
rect 6460 21904 6512 21913
rect 6644 21947 6696 21956
rect 6644 21913 6653 21947
rect 6653 21913 6687 21947
rect 6687 21913 6696 21947
rect 6644 21904 6696 21913
rect 16764 21947 16816 21956
rect 16764 21913 16773 21947
rect 16773 21913 16807 21947
rect 16807 21913 16816 21947
rect 16764 21904 16816 21913
rect 17224 22015 17276 22024
rect 17224 21981 17233 22015
rect 17233 21981 17267 22015
rect 17267 21981 17276 22015
rect 17224 21972 17276 21981
rect 17776 21972 17828 22024
rect 23664 22015 23716 22024
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 6828 21879 6880 21888
rect 6828 21845 6837 21879
rect 6837 21845 6871 21879
rect 6871 21845 6880 21879
rect 6828 21836 6880 21845
rect 11980 21836 12032 21888
rect 14188 21879 14240 21888
rect 14188 21845 14197 21879
rect 14197 21845 14231 21879
rect 14231 21845 14240 21879
rect 14188 21836 14240 21845
rect 14740 21836 14792 21888
rect 16672 21836 16724 21888
rect 23572 21836 23624 21888
rect 4473 21734 4525 21786
rect 4537 21734 4589 21786
rect 4601 21734 4653 21786
rect 4665 21734 4717 21786
rect 4729 21734 4781 21786
rect 10200 21734 10252 21786
rect 10264 21734 10316 21786
rect 10328 21734 10380 21786
rect 10392 21734 10444 21786
rect 10456 21734 10508 21786
rect 15927 21734 15979 21786
rect 15991 21734 16043 21786
rect 16055 21734 16107 21786
rect 16119 21734 16171 21786
rect 16183 21734 16235 21786
rect 21654 21734 21706 21786
rect 21718 21734 21770 21786
rect 21782 21734 21834 21786
rect 21846 21734 21898 21786
rect 21910 21734 21962 21786
rect 848 21496 900 21548
rect 9956 21564 10008 21616
rect 4528 21539 4580 21548
rect 4528 21505 4562 21539
rect 4562 21505 4580 21539
rect 4528 21496 4580 21505
rect 8944 21496 8996 21548
rect 9220 21496 9272 21548
rect 5540 21428 5592 21480
rect 6092 21428 6144 21480
rect 6644 21428 6696 21480
rect 11244 21428 11296 21480
rect 11980 21496 12032 21548
rect 15108 21564 15160 21616
rect 6000 21360 6052 21412
rect 6460 21360 6512 21412
rect 8944 21403 8996 21412
rect 8944 21369 8953 21403
rect 8953 21369 8987 21403
rect 8987 21369 8996 21403
rect 8944 21360 8996 21369
rect 12072 21403 12124 21412
rect 12072 21369 12081 21403
rect 12081 21369 12115 21403
rect 12115 21369 12124 21403
rect 15108 21428 15160 21480
rect 17408 21496 17460 21548
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 16764 21428 16816 21480
rect 17776 21428 17828 21480
rect 19892 21428 19944 21480
rect 23756 21496 23808 21548
rect 12072 21360 12124 21369
rect 14924 21360 14976 21412
rect 20720 21471 20772 21480
rect 20720 21437 20729 21471
rect 20729 21437 20763 21471
rect 20763 21437 20772 21471
rect 20720 21428 20772 21437
rect 20904 21471 20956 21480
rect 20904 21437 20913 21471
rect 20913 21437 20947 21471
rect 20947 21437 20956 21471
rect 20904 21428 20956 21437
rect 20812 21360 20864 21412
rect 4344 21335 4396 21344
rect 4344 21301 4353 21335
rect 4353 21301 4387 21335
rect 4387 21301 4396 21335
rect 4344 21292 4396 21301
rect 4436 21292 4488 21344
rect 7288 21292 7340 21344
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 10324 21292 10376 21344
rect 11796 21292 11848 21344
rect 11888 21292 11940 21344
rect 16948 21292 17000 21344
rect 19800 21292 19852 21344
rect 20536 21335 20588 21344
rect 20536 21301 20545 21335
rect 20545 21301 20579 21335
rect 20579 21301 20588 21335
rect 20536 21292 20588 21301
rect 23664 21335 23716 21344
rect 23664 21301 23673 21335
rect 23673 21301 23707 21335
rect 23707 21301 23716 21335
rect 23664 21292 23716 21301
rect 3813 21190 3865 21242
rect 3877 21190 3929 21242
rect 3941 21190 3993 21242
rect 4005 21190 4057 21242
rect 4069 21190 4121 21242
rect 9540 21190 9592 21242
rect 9604 21190 9656 21242
rect 9668 21190 9720 21242
rect 9732 21190 9784 21242
rect 9796 21190 9848 21242
rect 15267 21190 15319 21242
rect 15331 21190 15383 21242
rect 15395 21190 15447 21242
rect 15459 21190 15511 21242
rect 15523 21190 15575 21242
rect 20994 21190 21046 21242
rect 21058 21190 21110 21242
rect 21122 21190 21174 21242
rect 21186 21190 21238 21242
rect 21250 21190 21302 21242
rect 10324 21088 10376 21140
rect 15108 21131 15160 21140
rect 15108 21097 15117 21131
rect 15117 21097 15151 21131
rect 15151 21097 15160 21131
rect 15108 21088 15160 21097
rect 18052 21088 18104 21140
rect 4436 20995 4488 21004
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 5908 20952 5960 21004
rect 6092 20995 6144 21004
rect 6092 20961 6101 20995
rect 6101 20961 6135 20995
rect 6135 20961 6144 20995
rect 6092 20952 6144 20961
rect 6368 20995 6420 21004
rect 6368 20961 6377 20995
rect 6377 20961 6411 20995
rect 6411 20961 6420 20995
rect 6368 20952 6420 20961
rect 6828 20952 6880 21004
rect 7012 20995 7064 21004
rect 7012 20961 7021 20995
rect 7021 20961 7055 20995
rect 7055 20961 7064 20995
rect 7012 20952 7064 20961
rect 9220 20995 9272 21004
rect 9220 20961 9229 20995
rect 9229 20961 9263 20995
rect 9263 20961 9272 20995
rect 9220 20952 9272 20961
rect 9496 20995 9548 21004
rect 9496 20961 9505 20995
rect 9505 20961 9539 20995
rect 9539 20961 9548 20995
rect 9496 20952 9548 20961
rect 10692 20995 10744 21004
rect 10692 20961 10701 20995
rect 10701 20961 10735 20995
rect 10735 20961 10744 20995
rect 10692 20952 10744 20961
rect 11244 20995 11296 21004
rect 11244 20961 11253 20995
rect 11253 20961 11287 20995
rect 11287 20961 11296 20995
rect 11244 20952 11296 20961
rect 11888 20995 11940 21004
rect 11888 20961 11897 20995
rect 11897 20961 11931 20995
rect 11931 20961 11940 20995
rect 11888 20952 11940 20961
rect 12164 20952 12216 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 6000 20927 6052 20936
rect 6000 20893 6009 20927
rect 6009 20893 6043 20927
rect 6043 20893 6052 20927
rect 6000 20884 6052 20893
rect 7288 20927 7340 20936
rect 7288 20893 7297 20927
rect 7297 20893 7331 20927
rect 7331 20893 7340 20927
rect 7288 20884 7340 20893
rect 8944 20884 8996 20936
rect 10324 20927 10376 20936
rect 10324 20893 10333 20927
rect 10333 20893 10367 20927
rect 10367 20893 10376 20927
rect 10324 20884 10376 20893
rect 4528 20816 4580 20868
rect 7380 20816 7432 20868
rect 7472 20859 7524 20868
rect 7472 20825 7481 20859
rect 7481 20825 7515 20859
rect 7515 20825 7524 20859
rect 7472 20816 7524 20825
rect 11244 20816 11296 20868
rect 11796 20927 11848 20936
rect 11796 20893 11805 20927
rect 11805 20893 11839 20927
rect 11839 20893 11848 20927
rect 11796 20884 11848 20893
rect 3700 20748 3752 20800
rect 6736 20748 6788 20800
rect 11428 20791 11480 20800
rect 11428 20757 11437 20791
rect 11437 20757 11471 20791
rect 11471 20757 11480 20791
rect 11428 20748 11480 20757
rect 12072 20816 12124 20868
rect 14740 20995 14792 21004
rect 14740 20961 14749 20995
rect 14749 20961 14783 20995
rect 14783 20961 14792 20995
rect 14740 20952 14792 20961
rect 18144 21020 18196 21072
rect 17316 20995 17368 21004
rect 17316 20961 17325 20995
rect 17325 20961 17359 20995
rect 17359 20961 17368 20995
rect 17316 20952 17368 20961
rect 14648 20884 14700 20936
rect 15016 20884 15068 20936
rect 16948 20927 17000 20936
rect 16948 20893 16957 20927
rect 16957 20893 16991 20927
rect 16991 20893 17000 20927
rect 17592 20995 17644 21004
rect 17592 20961 17601 20995
rect 17601 20961 17635 20995
rect 17635 20961 17644 20995
rect 17592 20952 17644 20961
rect 20904 21020 20956 21072
rect 22744 20995 22796 21004
rect 22744 20961 22753 20995
rect 22753 20961 22787 20995
rect 22787 20961 22796 20995
rect 22744 20952 22796 20961
rect 16948 20884 17000 20893
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 20720 20884 20772 20936
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 23112 20927 23164 20936
rect 23112 20893 23120 20927
rect 23120 20893 23164 20927
rect 23112 20884 23164 20893
rect 23388 20884 23440 20936
rect 12624 20791 12676 20800
rect 12624 20757 12633 20791
rect 12633 20757 12667 20791
rect 12667 20757 12676 20791
rect 12624 20748 12676 20757
rect 13084 20791 13136 20800
rect 13084 20757 13093 20791
rect 13093 20757 13127 20791
rect 13127 20757 13136 20791
rect 13084 20748 13136 20757
rect 19432 20791 19484 20800
rect 19432 20757 19441 20791
rect 19441 20757 19475 20791
rect 19475 20757 19484 20791
rect 19432 20748 19484 20757
rect 19524 20748 19576 20800
rect 20720 20791 20772 20800
rect 20720 20757 20729 20791
rect 20729 20757 20763 20791
rect 20763 20757 20772 20791
rect 20720 20748 20772 20757
rect 21272 20748 21324 20800
rect 23480 20791 23532 20800
rect 23480 20757 23489 20791
rect 23489 20757 23523 20791
rect 23523 20757 23532 20791
rect 23480 20748 23532 20757
rect 4473 20646 4525 20698
rect 4537 20646 4589 20698
rect 4601 20646 4653 20698
rect 4665 20646 4717 20698
rect 4729 20646 4781 20698
rect 10200 20646 10252 20698
rect 10264 20646 10316 20698
rect 10328 20646 10380 20698
rect 10392 20646 10444 20698
rect 10456 20646 10508 20698
rect 15927 20646 15979 20698
rect 15991 20646 16043 20698
rect 16055 20646 16107 20698
rect 16119 20646 16171 20698
rect 16183 20646 16235 20698
rect 21654 20646 21706 20698
rect 21718 20646 21770 20698
rect 21782 20646 21834 20698
rect 21846 20646 21898 20698
rect 21910 20646 21962 20698
rect 7472 20544 7524 20596
rect 9496 20544 9548 20596
rect 14188 20587 14240 20596
rect 14188 20553 14197 20587
rect 14197 20553 14231 20587
rect 14231 20553 14240 20587
rect 14188 20544 14240 20553
rect 17316 20544 17368 20596
rect 19432 20587 19484 20596
rect 19432 20553 19441 20587
rect 19441 20553 19475 20587
rect 19475 20553 19484 20587
rect 19432 20544 19484 20553
rect 20720 20544 20772 20596
rect 3700 20408 3752 20460
rect 12624 20476 12676 20528
rect 19524 20476 19576 20528
rect 20536 20519 20588 20528
rect 20536 20485 20545 20519
rect 20545 20485 20579 20519
rect 20579 20485 20588 20519
rect 20536 20476 20588 20485
rect 6368 20408 6420 20460
rect 4344 20383 4396 20392
rect 4344 20349 4353 20383
rect 4353 20349 4387 20383
rect 4387 20349 4396 20383
rect 4344 20340 4396 20349
rect 9404 20383 9456 20392
rect 9404 20349 9413 20383
rect 9413 20349 9447 20383
rect 9447 20349 9456 20383
rect 9404 20340 9456 20349
rect 13084 20408 13136 20460
rect 14832 20408 14884 20460
rect 14924 20408 14976 20460
rect 20904 20476 20956 20528
rect 20812 20408 20864 20460
rect 6552 20315 6604 20324
rect 6552 20281 6561 20315
rect 6561 20281 6595 20315
rect 6595 20281 6604 20315
rect 6552 20272 6604 20281
rect 17500 20383 17552 20392
rect 17500 20349 17509 20383
rect 17509 20349 17543 20383
rect 17543 20349 17552 20383
rect 17500 20340 17552 20349
rect 17868 20340 17920 20392
rect 19800 20340 19852 20392
rect 19892 20383 19944 20392
rect 19892 20349 19901 20383
rect 19901 20349 19935 20383
rect 19935 20349 19944 20383
rect 19892 20340 19944 20349
rect 21272 20408 21324 20460
rect 3424 20247 3476 20256
rect 3424 20213 3433 20247
rect 3433 20213 3467 20247
rect 3467 20213 3476 20247
rect 3424 20204 3476 20213
rect 4252 20247 4304 20256
rect 4252 20213 4261 20247
rect 4261 20213 4295 20247
rect 4295 20213 4304 20247
rect 4252 20204 4304 20213
rect 4436 20204 4488 20256
rect 8944 20204 8996 20256
rect 10600 20247 10652 20256
rect 10600 20213 10609 20247
rect 10609 20213 10643 20247
rect 10643 20213 10652 20247
rect 10600 20204 10652 20213
rect 12716 20204 12768 20256
rect 14096 20204 14148 20256
rect 16764 20204 16816 20256
rect 18972 20247 19024 20256
rect 18972 20213 18981 20247
rect 18981 20213 19015 20247
rect 19015 20213 19024 20247
rect 18972 20204 19024 20213
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 3813 20102 3865 20154
rect 3877 20102 3929 20154
rect 3941 20102 3993 20154
rect 4005 20102 4057 20154
rect 4069 20102 4121 20154
rect 9540 20102 9592 20154
rect 9604 20102 9656 20154
rect 9668 20102 9720 20154
rect 9732 20102 9784 20154
rect 9796 20102 9848 20154
rect 15267 20102 15319 20154
rect 15331 20102 15383 20154
rect 15395 20102 15447 20154
rect 15459 20102 15511 20154
rect 15523 20102 15575 20154
rect 20994 20102 21046 20154
rect 21058 20102 21110 20154
rect 21122 20102 21174 20154
rect 21186 20102 21238 20154
rect 21250 20102 21302 20154
rect 14464 20000 14516 20052
rect 14924 20043 14976 20052
rect 14924 20009 14933 20043
rect 14933 20009 14967 20043
rect 14967 20009 14976 20043
rect 14924 20000 14976 20009
rect 16396 20000 16448 20052
rect 5356 19932 5408 19984
rect 9404 19932 9456 19984
rect 4252 19864 4304 19916
rect 848 19796 900 19848
rect 3424 19796 3476 19848
rect 4436 19839 4488 19848
rect 4436 19805 4445 19839
rect 4445 19805 4479 19839
rect 4479 19805 4488 19839
rect 4436 19796 4488 19805
rect 6368 19864 6420 19916
rect 6920 19907 6972 19916
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 8760 19864 8812 19916
rect 10600 19907 10652 19916
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 12164 19864 12216 19916
rect 14648 19907 14700 19916
rect 14648 19873 14657 19907
rect 14657 19873 14691 19907
rect 14691 19873 14700 19907
rect 14648 19864 14700 19873
rect 16764 19907 16816 19916
rect 16764 19873 16773 19907
rect 16773 19873 16807 19907
rect 16807 19873 16816 19907
rect 16764 19864 16816 19873
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 7104 19796 7156 19848
rect 11428 19796 11480 19848
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 14740 19796 14792 19848
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 16672 19839 16724 19848
rect 16672 19805 16681 19839
rect 16681 19805 16715 19839
rect 16715 19805 16724 19839
rect 16672 19796 16724 19805
rect 18788 19796 18840 19848
rect 4252 19728 4304 19780
rect 5080 19771 5132 19780
rect 5080 19737 5089 19771
rect 5089 19737 5123 19771
rect 5123 19737 5132 19771
rect 5080 19728 5132 19737
rect 10692 19728 10744 19780
rect 4804 19703 4856 19712
rect 4804 19669 4813 19703
rect 4813 19669 4847 19703
rect 4847 19669 4856 19703
rect 4804 19660 4856 19669
rect 9404 19660 9456 19712
rect 15844 19660 15896 19712
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 4473 19558 4525 19610
rect 4537 19558 4589 19610
rect 4601 19558 4653 19610
rect 4665 19558 4717 19610
rect 4729 19558 4781 19610
rect 10200 19558 10252 19610
rect 10264 19558 10316 19610
rect 10328 19558 10380 19610
rect 10392 19558 10444 19610
rect 10456 19558 10508 19610
rect 15927 19558 15979 19610
rect 15991 19558 16043 19610
rect 16055 19558 16107 19610
rect 16119 19558 16171 19610
rect 16183 19558 16235 19610
rect 21654 19558 21706 19610
rect 21718 19558 21770 19610
rect 21782 19558 21834 19610
rect 21846 19558 21898 19610
rect 21910 19558 21962 19610
rect 6920 19456 6972 19508
rect 7104 19499 7156 19508
rect 7104 19465 7113 19499
rect 7113 19465 7147 19499
rect 7147 19465 7156 19499
rect 7104 19456 7156 19465
rect 8944 19499 8996 19508
rect 8944 19465 8953 19499
rect 8953 19465 8987 19499
rect 8987 19465 8996 19499
rect 8944 19456 8996 19465
rect 9036 19499 9088 19508
rect 9036 19465 9045 19499
rect 9045 19465 9079 19499
rect 9079 19465 9088 19499
rect 9036 19456 9088 19465
rect 18788 19499 18840 19508
rect 18788 19465 18797 19499
rect 18797 19465 18831 19499
rect 18831 19465 18840 19499
rect 18788 19456 18840 19465
rect 23388 19499 23440 19508
rect 23388 19465 23397 19499
rect 23397 19465 23431 19499
rect 23431 19465 23440 19499
rect 23388 19456 23440 19465
rect 23664 19456 23716 19508
rect 7196 19388 7248 19440
rect 4344 19320 4396 19372
rect 14832 19320 14884 19372
rect 16948 19320 17000 19372
rect 18236 19320 18288 19372
rect 18972 19320 19024 19372
rect 23204 19363 23256 19372
rect 23204 19329 23213 19363
rect 23213 19329 23247 19363
rect 23247 19329 23256 19363
rect 23204 19320 23256 19329
rect 23296 19320 23348 19372
rect 3700 19295 3752 19304
rect 3700 19261 3709 19295
rect 3709 19261 3743 19295
rect 3743 19261 3752 19295
rect 3700 19252 3752 19261
rect 7012 19252 7064 19304
rect 8208 19252 8260 19304
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 1400 19159 1452 19168
rect 1400 19125 1409 19159
rect 1409 19125 1443 19159
rect 1443 19125 1452 19159
rect 1400 19116 1452 19125
rect 4160 19159 4212 19168
rect 4160 19125 4169 19159
rect 4169 19125 4203 19159
rect 4203 19125 4212 19159
rect 4160 19116 4212 19125
rect 6644 19159 6696 19168
rect 6644 19125 6653 19159
rect 6653 19125 6687 19159
rect 6687 19125 6696 19159
rect 6644 19116 6696 19125
rect 8944 19116 8996 19168
rect 3813 19014 3865 19066
rect 3877 19014 3929 19066
rect 3941 19014 3993 19066
rect 4005 19014 4057 19066
rect 4069 19014 4121 19066
rect 9540 19014 9592 19066
rect 9604 19014 9656 19066
rect 9668 19014 9720 19066
rect 9732 19014 9784 19066
rect 9796 19014 9848 19066
rect 15267 19014 15319 19066
rect 15331 19014 15383 19066
rect 15395 19014 15447 19066
rect 15459 19014 15511 19066
rect 15523 19014 15575 19066
rect 20994 19014 21046 19066
rect 21058 19014 21110 19066
rect 21122 19014 21174 19066
rect 21186 19014 21238 19066
rect 21250 19014 21302 19066
rect 5080 18912 5132 18964
rect 7196 18955 7248 18964
rect 7196 18921 7205 18955
rect 7205 18921 7239 18955
rect 7239 18921 7248 18955
rect 7196 18912 7248 18921
rect 9128 18955 9180 18964
rect 9128 18921 9137 18955
rect 9137 18921 9171 18955
rect 9171 18921 9180 18955
rect 9128 18912 9180 18921
rect 10048 18912 10100 18964
rect 15844 18912 15896 18964
rect 23204 18912 23256 18964
rect 4252 18776 4304 18828
rect 4436 18819 4488 18828
rect 4436 18785 4445 18819
rect 4445 18785 4479 18819
rect 4479 18785 4488 18819
rect 4436 18776 4488 18785
rect 4896 18776 4948 18828
rect 6644 18819 6696 18828
rect 6644 18785 6653 18819
rect 6653 18785 6687 18819
rect 6687 18785 6696 18819
rect 6644 18776 6696 18785
rect 12164 18819 12216 18828
rect 12164 18785 12173 18819
rect 12173 18785 12207 18819
rect 12207 18785 12216 18819
rect 12164 18776 12216 18785
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 4804 18708 4856 18760
rect 5080 18751 5132 18760
rect 5080 18717 5089 18751
rect 5089 18717 5123 18751
rect 5123 18717 5132 18751
rect 5080 18708 5132 18717
rect 6736 18751 6788 18760
rect 6736 18717 6745 18751
rect 6745 18717 6779 18751
rect 6779 18717 6788 18751
rect 6736 18708 6788 18717
rect 7012 18640 7064 18692
rect 8944 18751 8996 18760
rect 8944 18717 8953 18751
rect 8953 18717 8987 18751
rect 8987 18717 8996 18751
rect 8944 18708 8996 18717
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 12624 18819 12676 18828
rect 12624 18785 12633 18819
rect 12633 18785 12667 18819
rect 12667 18785 12676 18819
rect 12624 18776 12676 18785
rect 14096 18844 14148 18896
rect 14740 18844 14792 18896
rect 12716 18751 12768 18760
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 19800 18819 19852 18828
rect 19800 18785 19809 18819
rect 19809 18785 19843 18819
rect 19843 18785 19852 18819
rect 19800 18776 19852 18785
rect 12716 18708 12768 18717
rect 14096 18683 14148 18692
rect 14096 18649 14105 18683
rect 14105 18649 14139 18683
rect 14139 18649 14148 18683
rect 14096 18640 14148 18649
rect 14556 18640 14608 18692
rect 15292 18640 15344 18692
rect 18052 18708 18104 18760
rect 19248 18708 19300 18760
rect 23020 18776 23072 18828
rect 23204 18819 23256 18828
rect 23204 18785 23213 18819
rect 23213 18785 23247 18819
rect 23247 18785 23256 18819
rect 23204 18776 23256 18785
rect 19984 18708 20036 18760
rect 23480 18751 23532 18760
rect 23480 18717 23514 18751
rect 23514 18717 23532 18751
rect 23480 18708 23532 18717
rect 848 18572 900 18624
rect 4252 18572 4304 18624
rect 4988 18615 5040 18624
rect 4988 18581 4997 18615
rect 4997 18581 5031 18615
rect 5031 18581 5040 18615
rect 4988 18572 5040 18581
rect 7104 18615 7156 18624
rect 7104 18581 7113 18615
rect 7113 18581 7147 18615
rect 7147 18581 7156 18615
rect 7104 18572 7156 18581
rect 11520 18615 11572 18624
rect 11520 18581 11529 18615
rect 11529 18581 11563 18615
rect 11563 18581 11572 18615
rect 11520 18572 11572 18581
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 13268 18572 13320 18624
rect 14004 18572 14056 18624
rect 19524 18572 19576 18624
rect 22100 18640 22152 18692
rect 22376 18572 22428 18624
rect 22560 18615 22612 18624
rect 22560 18581 22569 18615
rect 22569 18581 22603 18615
rect 22603 18581 22612 18615
rect 22560 18572 22612 18581
rect 4473 18470 4525 18522
rect 4537 18470 4589 18522
rect 4601 18470 4653 18522
rect 4665 18470 4717 18522
rect 4729 18470 4781 18522
rect 10200 18470 10252 18522
rect 10264 18470 10316 18522
rect 10328 18470 10380 18522
rect 10392 18470 10444 18522
rect 10456 18470 10508 18522
rect 15927 18470 15979 18522
rect 15991 18470 16043 18522
rect 16055 18470 16107 18522
rect 16119 18470 16171 18522
rect 16183 18470 16235 18522
rect 21654 18470 21706 18522
rect 21718 18470 21770 18522
rect 21782 18470 21834 18522
rect 21846 18470 21898 18522
rect 21910 18470 21962 18522
rect 4252 18411 4304 18420
rect 4252 18377 4261 18411
rect 4261 18377 4295 18411
rect 4295 18377 4304 18411
rect 4252 18368 4304 18377
rect 5080 18368 5132 18420
rect 8668 18368 8720 18420
rect 14556 18411 14608 18420
rect 14556 18377 14565 18411
rect 14565 18377 14599 18411
rect 14599 18377 14608 18411
rect 14556 18368 14608 18377
rect 15292 18411 15344 18420
rect 15292 18377 15301 18411
rect 15301 18377 15335 18411
rect 15335 18377 15344 18411
rect 15292 18368 15344 18377
rect 18052 18368 18104 18420
rect 19524 18411 19576 18420
rect 19524 18377 19533 18411
rect 19533 18377 19567 18411
rect 19567 18377 19576 18411
rect 19524 18368 19576 18377
rect 19984 18411 20036 18420
rect 19984 18377 19993 18411
rect 19993 18377 20027 18411
rect 20027 18377 20036 18411
rect 19984 18368 20036 18377
rect 4344 18300 4396 18352
rect 9404 18300 9456 18352
rect 13268 18343 13320 18352
rect 13268 18309 13277 18343
rect 13277 18309 13311 18343
rect 13311 18309 13320 18343
rect 13268 18300 13320 18309
rect 3976 18164 4028 18216
rect 4988 18232 5040 18284
rect 11980 18232 12032 18284
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 5356 18164 5408 18216
rect 9404 18164 9456 18216
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 6092 18096 6144 18148
rect 8944 18096 8996 18148
rect 1400 18071 1452 18080
rect 1400 18037 1409 18071
rect 1409 18037 1443 18071
rect 1443 18037 1452 18071
rect 1400 18028 1452 18037
rect 13176 18028 13228 18080
rect 15844 18232 15896 18284
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 16948 18164 17000 18216
rect 15660 18139 15712 18148
rect 15660 18105 15669 18139
rect 15669 18105 15703 18139
rect 15703 18105 15712 18139
rect 15660 18096 15712 18105
rect 18144 18164 18196 18216
rect 19248 18164 19300 18216
rect 20904 18232 20956 18284
rect 22560 18232 22612 18284
rect 23572 18275 23624 18284
rect 23572 18241 23580 18275
rect 23580 18241 23624 18275
rect 23572 18232 23624 18241
rect 19800 18096 19852 18148
rect 22744 18164 22796 18216
rect 23112 18207 23164 18216
rect 23112 18173 23121 18207
rect 23121 18173 23155 18207
rect 23155 18173 23164 18207
rect 23112 18164 23164 18173
rect 22284 18096 22336 18148
rect 15844 18028 15896 18080
rect 16580 18028 16632 18080
rect 17868 18028 17920 18080
rect 21364 18071 21416 18080
rect 21364 18037 21373 18071
rect 21373 18037 21407 18071
rect 21407 18037 21416 18071
rect 21364 18028 21416 18037
rect 3813 17926 3865 17978
rect 3877 17926 3929 17978
rect 3941 17926 3993 17978
rect 4005 17926 4057 17978
rect 4069 17926 4121 17978
rect 9540 17926 9592 17978
rect 9604 17926 9656 17978
rect 9668 17926 9720 17978
rect 9732 17926 9784 17978
rect 9796 17926 9848 17978
rect 15267 17926 15319 17978
rect 15331 17926 15383 17978
rect 15395 17926 15447 17978
rect 15459 17926 15511 17978
rect 15523 17926 15575 17978
rect 20994 17926 21046 17978
rect 21058 17926 21110 17978
rect 21122 17926 21174 17978
rect 21186 17926 21238 17978
rect 21250 17926 21302 17978
rect 6092 17867 6144 17876
rect 6092 17833 6101 17867
rect 6101 17833 6135 17867
rect 6135 17833 6144 17867
rect 6092 17824 6144 17833
rect 7104 17824 7156 17876
rect 9864 17867 9916 17876
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 12624 17867 12676 17876
rect 12624 17833 12633 17867
rect 12633 17833 12667 17867
rect 12667 17833 12676 17867
rect 12624 17824 12676 17833
rect 13084 17867 13136 17876
rect 13084 17833 13093 17867
rect 13093 17833 13127 17867
rect 13127 17833 13136 17867
rect 13084 17824 13136 17833
rect 14740 17867 14792 17876
rect 14740 17833 14749 17867
rect 14749 17833 14783 17867
rect 14783 17833 14792 17867
rect 14740 17824 14792 17833
rect 17316 17824 17368 17876
rect 22100 17867 22152 17876
rect 22100 17833 22109 17867
rect 22109 17833 22143 17867
rect 22143 17833 22152 17867
rect 22100 17824 22152 17833
rect 22376 17824 22428 17876
rect 6828 17799 6880 17808
rect 6828 17765 6837 17799
rect 6837 17765 6871 17799
rect 6871 17765 6880 17799
rect 6828 17756 6880 17765
rect 8760 17756 8812 17808
rect 11060 17756 11112 17808
rect 6276 17663 6328 17672
rect 6276 17629 6285 17663
rect 6285 17629 6319 17663
rect 6319 17629 6328 17663
rect 6276 17620 6328 17629
rect 4804 17552 4856 17604
rect 8208 17731 8260 17740
rect 8208 17697 8217 17731
rect 8217 17697 8251 17731
rect 8251 17697 8260 17731
rect 8208 17688 8260 17697
rect 9404 17663 9456 17672
rect 9404 17629 9413 17663
rect 9413 17629 9447 17663
rect 9447 17629 9456 17663
rect 9404 17620 9456 17629
rect 11520 17620 11572 17672
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 12624 17620 12676 17672
rect 15200 17620 15252 17672
rect 18144 17756 18196 17808
rect 22192 17756 22244 17808
rect 22560 17756 22612 17808
rect 23664 17799 23716 17808
rect 23664 17765 23673 17799
rect 23673 17765 23707 17799
rect 23707 17765 23716 17799
rect 23664 17756 23716 17765
rect 16580 17688 16632 17740
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 17868 17663 17920 17672
rect 17868 17629 17877 17663
rect 17877 17629 17911 17663
rect 17911 17629 17920 17663
rect 17868 17620 17920 17629
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 6644 17484 6696 17493
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 12348 17552 12400 17604
rect 10784 17527 10836 17536
rect 10784 17493 10793 17527
rect 10793 17493 10827 17527
rect 10827 17493 10836 17527
rect 10784 17484 10836 17493
rect 4473 17382 4525 17434
rect 4537 17382 4589 17434
rect 4601 17382 4653 17434
rect 4665 17382 4717 17434
rect 4729 17382 4781 17434
rect 10200 17382 10252 17434
rect 10264 17382 10316 17434
rect 10328 17382 10380 17434
rect 10392 17382 10444 17434
rect 10456 17382 10508 17434
rect 15927 17382 15979 17434
rect 15991 17382 16043 17434
rect 16055 17382 16107 17434
rect 16119 17382 16171 17434
rect 16183 17382 16235 17434
rect 21654 17382 21706 17434
rect 21718 17382 21770 17434
rect 21782 17382 21834 17434
rect 21846 17382 21898 17434
rect 21910 17382 21962 17434
rect 6276 17280 6328 17332
rect 7012 17323 7064 17332
rect 7012 17289 7021 17323
rect 7021 17289 7055 17323
rect 7055 17289 7064 17323
rect 7012 17280 7064 17289
rect 10784 17280 10836 17332
rect 15200 17280 15252 17332
rect 6644 17212 6696 17264
rect 13544 17212 13596 17264
rect 23572 17280 23624 17332
rect 848 17144 900 17196
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 6828 17144 6880 17196
rect 12624 17187 12676 17196
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 12716 17144 12768 17196
rect 13636 17144 13688 17196
rect 17868 17212 17920 17264
rect 18236 17144 18288 17196
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 4804 17119 4856 17128
rect 4804 17085 4813 17119
rect 4813 17085 4847 17119
rect 4847 17085 4856 17119
rect 4804 17076 4856 17085
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 12072 17119 12124 17128
rect 12072 17085 12081 17119
rect 12081 17085 12115 17119
rect 12115 17085 12124 17119
rect 12072 17076 12124 17085
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 13728 17076 13780 17128
rect 16212 17076 16264 17128
rect 11796 17008 11848 17060
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 11060 16940 11112 16992
rect 12348 17008 12400 17060
rect 16120 17008 16172 17060
rect 19524 17144 19576 17196
rect 12900 16940 12952 16992
rect 15936 16940 15988 16992
rect 18236 16940 18288 16992
rect 23664 17051 23716 17060
rect 23664 17017 23673 17051
rect 23673 17017 23707 17051
rect 23707 17017 23716 17051
rect 23664 17008 23716 17017
rect 23848 16940 23900 16992
rect 3813 16838 3865 16890
rect 3877 16838 3929 16890
rect 3941 16838 3993 16890
rect 4005 16838 4057 16890
rect 4069 16838 4121 16890
rect 9540 16838 9592 16890
rect 9604 16838 9656 16890
rect 9668 16838 9720 16890
rect 9732 16838 9784 16890
rect 9796 16838 9848 16890
rect 15267 16838 15319 16890
rect 15331 16838 15383 16890
rect 15395 16838 15447 16890
rect 15459 16838 15511 16890
rect 15523 16838 15575 16890
rect 20994 16838 21046 16890
rect 21058 16838 21110 16890
rect 21122 16838 21174 16890
rect 21186 16838 21238 16890
rect 21250 16838 21302 16890
rect 4896 16736 4948 16788
rect 7196 16736 7248 16788
rect 9404 16779 9456 16788
rect 9404 16745 9413 16779
rect 9413 16745 9447 16779
rect 9447 16745 9456 16779
rect 9404 16736 9456 16745
rect 12072 16736 12124 16788
rect 5448 16668 5500 16720
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 8208 16668 8260 16720
rect 11060 16668 11112 16720
rect 5356 16600 5408 16609
rect 8852 16600 8904 16652
rect 848 16532 900 16584
rect 9772 16507 9824 16516
rect 9772 16473 9781 16507
rect 9781 16473 9815 16507
rect 9815 16473 9824 16507
rect 9772 16464 9824 16473
rect 5172 16439 5224 16448
rect 5172 16405 5181 16439
rect 5181 16405 5215 16439
rect 5215 16405 5224 16439
rect 5172 16396 5224 16405
rect 6920 16396 6972 16448
rect 7564 16439 7616 16448
rect 7564 16405 7573 16439
rect 7573 16405 7607 16439
rect 7607 16405 7616 16439
rect 7564 16396 7616 16405
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 9864 16396 9916 16405
rect 10048 16532 10100 16584
rect 12348 16575 12400 16584
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 12348 16532 12400 16541
rect 12624 16736 12676 16788
rect 15844 16736 15896 16788
rect 18328 16736 18380 16788
rect 19524 16779 19576 16788
rect 19524 16745 19533 16779
rect 19533 16745 19567 16779
rect 19567 16745 19576 16779
rect 19524 16736 19576 16745
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 15936 16643 15988 16652
rect 15936 16609 15945 16643
rect 15945 16609 15979 16643
rect 15979 16609 15988 16643
rect 15936 16600 15988 16609
rect 16212 16668 16264 16720
rect 22008 16668 22060 16720
rect 18328 16600 18380 16652
rect 19800 16600 19852 16652
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 16120 16532 16172 16584
rect 18420 16532 18472 16584
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 20720 16575 20772 16584
rect 20720 16541 20729 16575
rect 20729 16541 20763 16575
rect 20763 16541 20772 16575
rect 20720 16532 20772 16541
rect 23664 16575 23716 16584
rect 23664 16541 23673 16575
rect 23673 16541 23707 16575
rect 23707 16541 23716 16575
rect 23664 16532 23716 16541
rect 11888 16396 11940 16448
rect 17960 16439 18012 16448
rect 17960 16405 17969 16439
rect 17969 16405 18003 16439
rect 18003 16405 18012 16439
rect 17960 16396 18012 16405
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 23756 16464 23808 16516
rect 19892 16439 19944 16448
rect 19892 16405 19901 16439
rect 19901 16405 19935 16439
rect 19935 16405 19944 16439
rect 19892 16396 19944 16405
rect 19984 16439 20036 16448
rect 19984 16405 19993 16439
rect 19993 16405 20027 16439
rect 20027 16405 20036 16439
rect 19984 16396 20036 16405
rect 23480 16439 23532 16448
rect 23480 16405 23489 16439
rect 23489 16405 23523 16439
rect 23523 16405 23532 16439
rect 23480 16396 23532 16405
rect 4473 16294 4525 16346
rect 4537 16294 4589 16346
rect 4601 16294 4653 16346
rect 4665 16294 4717 16346
rect 4729 16294 4781 16346
rect 10200 16294 10252 16346
rect 10264 16294 10316 16346
rect 10328 16294 10380 16346
rect 10392 16294 10444 16346
rect 10456 16294 10508 16346
rect 15927 16294 15979 16346
rect 15991 16294 16043 16346
rect 16055 16294 16107 16346
rect 16119 16294 16171 16346
rect 16183 16294 16235 16346
rect 21654 16294 21706 16346
rect 21718 16294 21770 16346
rect 21782 16294 21834 16346
rect 21846 16294 21898 16346
rect 21910 16294 21962 16346
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 7564 16192 7616 16244
rect 9864 16192 9916 16244
rect 10048 16192 10100 16244
rect 12348 16235 12400 16244
rect 12348 16201 12357 16235
rect 12357 16201 12391 16235
rect 12391 16201 12400 16235
rect 12348 16192 12400 16201
rect 12716 16235 12768 16244
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 12900 16192 12952 16244
rect 15752 16192 15804 16244
rect 17960 16192 18012 16244
rect 18788 16192 18840 16244
rect 19984 16192 20036 16244
rect 20720 16192 20772 16244
rect 5080 16124 5132 16176
rect 848 16056 900 16108
rect 3240 16056 3292 16108
rect 5448 16056 5500 16108
rect 6828 16056 6880 16108
rect 4252 15988 4304 16040
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 7288 16056 7340 16108
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 14096 16099 14148 16108
rect 14096 16065 14105 16099
rect 14105 16065 14139 16099
rect 14139 16065 14148 16099
rect 14096 16056 14148 16065
rect 18512 16099 18564 16108
rect 18512 16065 18521 16099
rect 18521 16065 18555 16099
rect 18555 16065 18564 16099
rect 18512 16056 18564 16065
rect 11060 15988 11112 16040
rect 12992 16031 13044 16040
rect 12992 15997 13001 16031
rect 13001 15997 13035 16031
rect 13035 15997 13044 16031
rect 12992 15988 13044 15997
rect 13728 15988 13780 16040
rect 17960 15988 18012 16040
rect 18144 15988 18196 16040
rect 19064 15988 19116 16040
rect 21548 15988 21600 16040
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22192 16056 22244 16065
rect 23664 16099 23716 16108
rect 23664 16065 23673 16099
rect 23673 16065 23707 16099
rect 23707 16065 23716 16099
rect 23664 16056 23716 16065
rect 22008 15988 22060 16040
rect 7380 15920 7432 15972
rect 6460 15852 6512 15904
rect 23572 15852 23624 15904
rect 3813 15750 3865 15802
rect 3877 15750 3929 15802
rect 3941 15750 3993 15802
rect 4005 15750 4057 15802
rect 4069 15750 4121 15802
rect 9540 15750 9592 15802
rect 9604 15750 9656 15802
rect 9668 15750 9720 15802
rect 9732 15750 9784 15802
rect 9796 15750 9848 15802
rect 15267 15750 15319 15802
rect 15331 15750 15383 15802
rect 15395 15750 15447 15802
rect 15459 15750 15511 15802
rect 15523 15750 15575 15802
rect 20994 15750 21046 15802
rect 21058 15750 21110 15802
rect 21122 15750 21174 15802
rect 21186 15750 21238 15802
rect 21250 15750 21302 15802
rect 3240 15691 3292 15700
rect 3240 15657 3249 15691
rect 3249 15657 3283 15691
rect 3283 15657 3292 15691
rect 3240 15648 3292 15657
rect 4988 15691 5040 15700
rect 4988 15657 4997 15691
rect 4997 15657 5031 15691
rect 5031 15657 5040 15691
rect 4988 15648 5040 15657
rect 5080 15691 5132 15700
rect 5080 15657 5089 15691
rect 5089 15657 5123 15691
rect 5123 15657 5132 15691
rect 5080 15648 5132 15657
rect 5448 15623 5500 15632
rect 5448 15589 5457 15623
rect 5457 15589 5491 15623
rect 5491 15589 5500 15623
rect 5448 15580 5500 15589
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 6920 15648 6972 15657
rect 8024 15648 8076 15700
rect 9864 15648 9916 15700
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 19892 15648 19944 15700
rect 7012 15580 7064 15632
rect 22192 15623 22244 15632
rect 22192 15589 22201 15623
rect 22201 15589 22235 15623
rect 22235 15589 22244 15623
rect 22192 15580 22244 15589
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 3424 15487 3476 15496
rect 3424 15453 3433 15487
rect 3433 15453 3467 15487
rect 3467 15453 3476 15487
rect 3424 15444 3476 15453
rect 5356 15512 5408 15564
rect 6644 15512 6696 15564
rect 7288 15555 7340 15564
rect 7288 15521 7297 15555
rect 7297 15521 7331 15555
rect 7331 15521 7340 15555
rect 7288 15512 7340 15521
rect 8760 15555 8812 15564
rect 8760 15521 8769 15555
rect 8769 15521 8803 15555
rect 8803 15521 8812 15555
rect 8760 15512 8812 15521
rect 11060 15512 11112 15564
rect 14832 15512 14884 15564
rect 15660 15512 15712 15564
rect 18880 15512 18932 15564
rect 21548 15555 21600 15564
rect 21548 15521 21557 15555
rect 21557 15521 21591 15555
rect 21591 15521 21600 15555
rect 21548 15512 21600 15521
rect 4252 15444 4304 15496
rect 3608 15376 3660 15428
rect 3424 15308 3476 15360
rect 6460 15419 6512 15428
rect 6460 15385 6469 15419
rect 6469 15385 6503 15419
rect 6503 15385 6512 15419
rect 6460 15376 6512 15385
rect 6828 15444 6880 15496
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 17960 15444 18012 15453
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 23388 15444 23440 15496
rect 10692 15376 10744 15428
rect 4804 15308 4856 15360
rect 10600 15308 10652 15360
rect 14464 15351 14516 15360
rect 14464 15317 14473 15351
rect 14473 15317 14507 15351
rect 14507 15317 14516 15351
rect 14464 15308 14516 15317
rect 15200 15308 15252 15360
rect 17132 15308 17184 15360
rect 21364 15351 21416 15360
rect 21364 15317 21373 15351
rect 21373 15317 21407 15351
rect 21407 15317 21416 15351
rect 21364 15308 21416 15317
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 21548 15308 21600 15360
rect 23664 15308 23716 15360
rect 4473 15206 4525 15258
rect 4537 15206 4589 15258
rect 4601 15206 4653 15258
rect 4665 15206 4717 15258
rect 4729 15206 4781 15258
rect 10200 15206 10252 15258
rect 10264 15206 10316 15258
rect 10328 15206 10380 15258
rect 10392 15206 10444 15258
rect 10456 15206 10508 15258
rect 15927 15206 15979 15258
rect 15991 15206 16043 15258
rect 16055 15206 16107 15258
rect 16119 15206 16171 15258
rect 16183 15206 16235 15258
rect 21654 15206 21706 15258
rect 21718 15206 21770 15258
rect 21782 15206 21834 15258
rect 21846 15206 21898 15258
rect 21910 15206 21962 15258
rect 4804 15104 4856 15156
rect 7288 15104 7340 15156
rect 7380 15147 7432 15156
rect 7380 15113 7389 15147
rect 7389 15113 7423 15147
rect 7423 15113 7432 15147
rect 7380 15104 7432 15113
rect 8760 15104 8812 15156
rect 10600 15147 10652 15156
rect 10600 15113 10609 15147
rect 10609 15113 10643 15147
rect 10643 15113 10652 15147
rect 10600 15104 10652 15113
rect 10692 15147 10744 15156
rect 10692 15113 10701 15147
rect 10701 15113 10735 15147
rect 10735 15113 10744 15147
rect 10692 15104 10744 15113
rect 18052 15104 18104 15156
rect 21364 15104 21416 15156
rect 3608 14968 3660 15020
rect 3424 14900 3476 14952
rect 3700 14900 3752 14952
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 5264 14968 5316 15020
rect 8668 15036 8720 15088
rect 12440 15036 12492 15088
rect 13084 15036 13136 15088
rect 17960 15036 18012 15088
rect 7472 14943 7524 14952
rect 7472 14909 7481 14943
rect 7481 14909 7515 14943
rect 7515 14909 7524 14943
rect 7472 14900 7524 14909
rect 9404 14968 9456 15020
rect 11888 15011 11940 15020
rect 11888 14977 11932 15011
rect 11932 14977 11940 15011
rect 11888 14968 11940 14977
rect 15660 14968 15712 15020
rect 10876 14943 10928 14952
rect 10876 14909 10885 14943
rect 10885 14909 10919 14943
rect 10919 14909 10928 14943
rect 10876 14900 10928 14909
rect 17868 14968 17920 15020
rect 18052 15011 18104 15020
rect 18052 14977 18061 15011
rect 18061 14977 18095 15011
rect 18095 14977 18104 15011
rect 18052 14968 18104 14977
rect 10232 14832 10284 14884
rect 12348 14832 12400 14884
rect 17592 14832 17644 14884
rect 18420 14900 18472 14952
rect 18512 14943 18564 14952
rect 18512 14909 18521 14943
rect 18521 14909 18555 14943
rect 18555 14909 18564 14943
rect 18512 14900 18564 14909
rect 21548 15036 21600 15088
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 21640 15011 21692 15020
rect 21640 14977 21649 15011
rect 21649 14977 21683 15011
rect 21683 14977 21692 15011
rect 21640 14968 21692 14977
rect 23572 15011 23624 15020
rect 23572 14977 23580 15011
rect 23580 14977 23624 15011
rect 22008 14900 22060 14952
rect 22100 14943 22152 14952
rect 22100 14909 22109 14943
rect 22109 14909 22143 14943
rect 22143 14909 22152 14943
rect 22100 14900 22152 14909
rect 17868 14832 17920 14884
rect 23572 14968 23624 14977
rect 23296 14900 23348 14952
rect 10876 14764 10928 14816
rect 12808 14764 12860 14816
rect 17316 14764 17368 14816
rect 22284 14764 22336 14816
rect 3813 14662 3865 14714
rect 3877 14662 3929 14714
rect 3941 14662 3993 14714
rect 4005 14662 4057 14714
rect 4069 14662 4121 14714
rect 9540 14662 9592 14714
rect 9604 14662 9656 14714
rect 9668 14662 9720 14714
rect 9732 14662 9784 14714
rect 9796 14662 9848 14714
rect 15267 14662 15319 14714
rect 15331 14662 15383 14714
rect 15395 14662 15447 14714
rect 15459 14662 15511 14714
rect 15523 14662 15575 14714
rect 20994 14662 21046 14714
rect 21058 14662 21110 14714
rect 21122 14662 21174 14714
rect 21186 14662 21238 14714
rect 21250 14662 21302 14714
rect 3608 14603 3660 14612
rect 3608 14569 3617 14603
rect 3617 14569 3651 14603
rect 3651 14569 3660 14603
rect 3608 14560 3660 14569
rect 3700 14560 3752 14612
rect 6644 14603 6696 14612
rect 6644 14569 6653 14603
rect 6653 14569 6687 14603
rect 6687 14569 6696 14603
rect 6644 14560 6696 14569
rect 7472 14560 7524 14612
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 10048 14560 10100 14612
rect 10876 14560 10928 14612
rect 12348 14603 12400 14612
rect 12348 14569 12357 14603
rect 12357 14569 12391 14603
rect 12391 14569 12400 14603
rect 12348 14560 12400 14569
rect 14464 14560 14516 14612
rect 15108 14603 15160 14612
rect 15108 14569 15117 14603
rect 15117 14569 15151 14603
rect 15151 14569 15160 14603
rect 15108 14560 15160 14569
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 18420 14603 18472 14612
rect 18420 14569 18429 14603
rect 18429 14569 18463 14603
rect 18463 14569 18472 14603
rect 18420 14560 18472 14569
rect 21456 14603 21508 14612
rect 21456 14569 21465 14603
rect 21465 14569 21499 14603
rect 21499 14569 21508 14603
rect 21456 14560 21508 14569
rect 21640 14560 21692 14612
rect 5080 14424 5132 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 9956 14424 10008 14476
rect 10692 14424 10744 14476
rect 11060 14492 11112 14544
rect 12440 14424 12492 14476
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 12992 14467 13044 14476
rect 12992 14433 13001 14467
rect 13001 14433 13035 14467
rect 13035 14433 13044 14467
rect 12992 14424 13044 14433
rect 15660 14492 15712 14544
rect 23664 14560 23716 14612
rect 15568 14467 15620 14476
rect 15568 14433 15577 14467
rect 15577 14433 15611 14467
rect 15611 14433 15620 14467
rect 15568 14424 15620 14433
rect 848 14356 900 14408
rect 4344 14220 4396 14272
rect 7012 14399 7064 14408
rect 7012 14365 7021 14399
rect 7021 14365 7055 14399
rect 7055 14365 7064 14399
rect 7012 14356 7064 14365
rect 7380 14356 7432 14408
rect 10232 14399 10284 14408
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 9956 14288 10008 14340
rect 11888 14356 11940 14408
rect 13820 14356 13872 14408
rect 15660 14356 15712 14408
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 17592 14399 17644 14408
rect 17592 14365 17601 14399
rect 17601 14365 17635 14399
rect 17635 14365 17644 14399
rect 17592 14356 17644 14365
rect 14096 14288 14148 14340
rect 22284 14535 22336 14544
rect 22284 14501 22293 14535
rect 22293 14501 22327 14535
rect 22327 14501 22336 14535
rect 22284 14492 22336 14501
rect 23112 14467 23164 14476
rect 11796 14220 11848 14272
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14464 14220 14516 14229
rect 17868 14220 17920 14272
rect 22100 14399 22152 14408
rect 22100 14365 22109 14399
rect 22109 14365 22143 14399
rect 22143 14365 22152 14399
rect 22100 14356 22152 14365
rect 22192 14356 22244 14408
rect 23112 14433 23121 14467
rect 23121 14433 23155 14467
rect 23155 14433 23164 14467
rect 23112 14424 23164 14433
rect 23480 14399 23532 14408
rect 23480 14365 23514 14399
rect 23514 14365 23532 14399
rect 23480 14356 23532 14365
rect 22192 14220 22244 14272
rect 4473 14118 4525 14170
rect 4537 14118 4589 14170
rect 4601 14118 4653 14170
rect 4665 14118 4717 14170
rect 4729 14118 4781 14170
rect 10200 14118 10252 14170
rect 10264 14118 10316 14170
rect 10328 14118 10380 14170
rect 10392 14118 10444 14170
rect 10456 14118 10508 14170
rect 15927 14118 15979 14170
rect 15991 14118 16043 14170
rect 16055 14118 16107 14170
rect 16119 14118 16171 14170
rect 16183 14118 16235 14170
rect 21654 14118 21706 14170
rect 21718 14118 21770 14170
rect 21782 14118 21834 14170
rect 21846 14118 21898 14170
rect 21910 14118 21962 14170
rect 4344 14016 4396 14068
rect 11980 14016 12032 14068
rect 14464 14016 14516 14068
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 11796 13880 11848 13932
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14096 13812 14148 13864
rect 15568 13880 15620 13932
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 7196 13744 7248 13796
rect 12992 13744 13044 13796
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 17868 13923 17920 13932
rect 17868 13889 17877 13923
rect 17877 13889 17911 13923
rect 17911 13889 17920 13923
rect 17868 13880 17920 13889
rect 23388 13923 23440 13932
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 23664 13923 23716 13932
rect 23664 13889 23673 13923
rect 23673 13889 23707 13923
rect 23707 13889 23716 13923
rect 23664 13880 23716 13889
rect 17224 13744 17276 13796
rect 15752 13676 15804 13728
rect 17040 13676 17092 13728
rect 23204 13719 23256 13728
rect 23204 13685 23213 13719
rect 23213 13685 23247 13719
rect 23247 13685 23256 13719
rect 23204 13676 23256 13685
rect 3813 13574 3865 13626
rect 3877 13574 3929 13626
rect 3941 13574 3993 13626
rect 4005 13574 4057 13626
rect 4069 13574 4121 13626
rect 9540 13574 9592 13626
rect 9604 13574 9656 13626
rect 9668 13574 9720 13626
rect 9732 13574 9784 13626
rect 9796 13574 9848 13626
rect 15267 13574 15319 13626
rect 15331 13574 15383 13626
rect 15395 13574 15447 13626
rect 15459 13574 15511 13626
rect 15523 13574 15575 13626
rect 20994 13574 21046 13626
rect 21058 13574 21110 13626
rect 21122 13574 21174 13626
rect 21186 13574 21238 13626
rect 21250 13574 21302 13626
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 17132 13472 17184 13524
rect 12992 13336 13044 13388
rect 13268 13336 13320 13388
rect 14096 13336 14148 13388
rect 848 13268 900 13320
rect 7012 13311 7064 13320
rect 7012 13277 7030 13311
rect 7030 13277 7064 13311
rect 7012 13268 7064 13277
rect 23204 13404 23256 13456
rect 19984 13336 20036 13388
rect 15752 13268 15804 13320
rect 17224 13311 17276 13320
rect 17224 13277 17258 13311
rect 17258 13277 17276 13311
rect 17224 13268 17276 13277
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 20628 13268 20680 13320
rect 23664 13311 23716 13320
rect 23664 13277 23673 13311
rect 23673 13277 23707 13311
rect 23707 13277 23716 13311
rect 23664 13268 23716 13277
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 6920 13132 6972 13184
rect 15844 13132 15896 13184
rect 19156 13132 19208 13184
rect 20720 13132 20772 13184
rect 4473 13030 4525 13082
rect 4537 13030 4589 13082
rect 4601 13030 4653 13082
rect 4665 13030 4717 13082
rect 4729 13030 4781 13082
rect 10200 13030 10252 13082
rect 10264 13030 10316 13082
rect 10328 13030 10380 13082
rect 10392 13030 10444 13082
rect 10456 13030 10508 13082
rect 15927 13030 15979 13082
rect 15991 13030 16043 13082
rect 16055 13030 16107 13082
rect 16119 13030 16171 13082
rect 16183 13030 16235 13082
rect 21654 13030 21706 13082
rect 21718 13030 21770 13082
rect 21782 13030 21834 13082
rect 21846 13030 21898 13082
rect 21910 13030 21962 13082
rect 1584 12860 1636 12912
rect 6920 12971 6972 12980
rect 6920 12937 6929 12971
rect 6929 12937 6963 12971
rect 6963 12937 6972 12971
rect 6920 12928 6972 12937
rect 9956 12928 10008 12980
rect 14096 12928 14148 12980
rect 19156 12971 19208 12980
rect 19156 12937 19165 12971
rect 19165 12937 19199 12971
rect 19199 12937 19208 12971
rect 19156 12928 19208 12937
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 4804 12792 4856 12844
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 19432 12860 19484 12912
rect 19984 12903 20036 12912
rect 19984 12869 19993 12903
rect 19993 12869 20027 12903
rect 20027 12869 20036 12903
rect 20628 12971 20680 12980
rect 20628 12937 20637 12971
rect 20637 12937 20671 12971
rect 20671 12937 20680 12971
rect 20628 12928 20680 12937
rect 20720 12971 20772 12980
rect 20720 12937 20729 12971
rect 20729 12937 20763 12971
rect 20763 12937 20772 12971
rect 20720 12928 20772 12937
rect 19984 12860 20036 12869
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 10876 12792 10928 12844
rect 14924 12792 14976 12844
rect 21364 12792 21416 12844
rect 4712 12656 4764 12708
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 6920 12724 6972 12776
rect 7104 12724 7156 12776
rect 7380 12699 7432 12708
rect 7380 12665 7389 12699
rect 7389 12665 7423 12699
rect 7423 12665 7432 12699
rect 7380 12656 7432 12665
rect 4344 12588 4396 12640
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 19064 12724 19116 12776
rect 23388 12792 23440 12844
rect 8300 12656 8352 12708
rect 17040 12656 17092 12708
rect 23204 12656 23256 12708
rect 8208 12588 8260 12640
rect 11060 12588 11112 12640
rect 18236 12588 18288 12640
rect 20904 12588 20956 12640
rect 3813 12486 3865 12538
rect 3877 12486 3929 12538
rect 3941 12486 3993 12538
rect 4005 12486 4057 12538
rect 4069 12486 4121 12538
rect 9540 12486 9592 12538
rect 9604 12486 9656 12538
rect 9668 12486 9720 12538
rect 9732 12486 9784 12538
rect 9796 12486 9848 12538
rect 15267 12486 15319 12538
rect 15331 12486 15383 12538
rect 15395 12486 15447 12538
rect 15459 12486 15511 12538
rect 15523 12486 15575 12538
rect 20994 12486 21046 12538
rect 21058 12486 21110 12538
rect 21122 12486 21174 12538
rect 21186 12486 21238 12538
rect 21250 12486 21302 12538
rect 5356 12384 5408 12436
rect 6920 12384 6972 12436
rect 7288 12384 7340 12436
rect 10416 12384 10468 12436
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 7380 12316 7432 12368
rect 8208 12248 8260 12300
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 5540 12044 5592 12096
rect 8484 12155 8536 12164
rect 8484 12121 8493 12155
rect 8493 12121 8527 12155
rect 8527 12121 8536 12155
rect 8484 12112 8536 12121
rect 10048 12112 10100 12164
rect 10600 12180 10652 12232
rect 11612 12155 11664 12164
rect 11612 12121 11621 12155
rect 11621 12121 11655 12155
rect 11655 12121 11664 12155
rect 11612 12112 11664 12121
rect 15568 12248 15620 12300
rect 16488 12248 16540 12300
rect 18972 12248 19024 12300
rect 19432 12248 19484 12300
rect 12624 12180 12676 12232
rect 15752 12180 15804 12232
rect 17040 12180 17092 12232
rect 11888 12112 11940 12164
rect 19984 12316 20036 12368
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 22192 12248 22244 12300
rect 21364 12180 21416 12232
rect 7380 12087 7432 12096
rect 7380 12053 7389 12087
rect 7389 12053 7423 12087
rect 7423 12053 7432 12087
rect 7380 12044 7432 12053
rect 11428 12087 11480 12096
rect 11428 12053 11437 12087
rect 11437 12053 11471 12087
rect 11471 12053 11480 12087
rect 11428 12044 11480 12053
rect 12440 12044 12492 12096
rect 17132 12044 17184 12096
rect 20168 12044 20220 12096
rect 4473 11942 4525 11994
rect 4537 11942 4589 11994
rect 4601 11942 4653 11994
rect 4665 11942 4717 11994
rect 4729 11942 4781 11994
rect 10200 11942 10252 11994
rect 10264 11942 10316 11994
rect 10328 11942 10380 11994
rect 10392 11942 10444 11994
rect 10456 11942 10508 11994
rect 15927 11942 15979 11994
rect 15991 11942 16043 11994
rect 16055 11942 16107 11994
rect 16119 11942 16171 11994
rect 16183 11942 16235 11994
rect 21654 11942 21706 11994
rect 21718 11942 21770 11994
rect 21782 11942 21834 11994
rect 21846 11942 21898 11994
rect 21910 11942 21962 11994
rect 4804 11840 4856 11892
rect 8484 11840 8536 11892
rect 10048 11840 10100 11892
rect 10600 11840 10652 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 12808 11840 12860 11892
rect 13820 11840 13872 11892
rect 5448 11772 5500 11824
rect 8208 11772 8260 11824
rect 848 11704 900 11756
rect 4160 11704 4212 11756
rect 4344 11704 4396 11756
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 5448 11636 5500 11688
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 7104 11636 7156 11688
rect 7748 11568 7800 11620
rect 4620 11500 4672 11552
rect 4988 11500 5040 11552
rect 5816 11500 5868 11552
rect 7656 11500 7708 11552
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 11612 11636 11664 11688
rect 11888 11611 11940 11620
rect 11888 11577 11897 11611
rect 11897 11577 11931 11611
rect 11931 11577 11940 11611
rect 11888 11568 11940 11577
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 15752 11704 15804 11756
rect 13084 11568 13136 11620
rect 16028 11611 16080 11620
rect 16028 11577 16037 11611
rect 16037 11577 16071 11611
rect 16071 11577 16080 11611
rect 16028 11568 16080 11577
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 17040 11815 17092 11824
rect 17040 11781 17049 11815
rect 17049 11781 17083 11815
rect 17083 11781 17092 11815
rect 17040 11772 17092 11781
rect 20168 11815 20220 11824
rect 20168 11781 20177 11815
rect 20177 11781 20211 11815
rect 20211 11781 20220 11815
rect 20168 11772 20220 11781
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 23664 11747 23716 11756
rect 23664 11713 23673 11747
rect 23673 11713 23707 11747
rect 23707 11713 23716 11747
rect 23664 11704 23716 11713
rect 18512 11568 18564 11620
rect 10048 11500 10100 11552
rect 11520 11543 11572 11552
rect 11520 11509 11529 11543
rect 11529 11509 11563 11543
rect 11563 11509 11572 11543
rect 11520 11500 11572 11509
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 18420 11500 18472 11552
rect 20720 11500 20772 11552
rect 3813 11398 3865 11450
rect 3877 11398 3929 11450
rect 3941 11398 3993 11450
rect 4005 11398 4057 11450
rect 4069 11398 4121 11450
rect 9540 11398 9592 11450
rect 9604 11398 9656 11450
rect 9668 11398 9720 11450
rect 9732 11398 9784 11450
rect 9796 11398 9848 11450
rect 15267 11398 15319 11450
rect 15331 11398 15383 11450
rect 15395 11398 15447 11450
rect 15459 11398 15511 11450
rect 15523 11398 15575 11450
rect 20994 11398 21046 11450
rect 21058 11398 21110 11450
rect 21122 11398 21174 11450
rect 21186 11398 21238 11450
rect 21250 11398 21302 11450
rect 4896 11296 4948 11348
rect 10508 11296 10560 11348
rect 11060 11296 11112 11348
rect 9312 11228 9364 11280
rect 4344 11160 4396 11212
rect 5080 11203 5132 11212
rect 5080 11169 5089 11203
rect 5089 11169 5123 11203
rect 5123 11169 5132 11203
rect 5080 11160 5132 11169
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 4620 11092 4672 11144
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 7656 11203 7708 11212
rect 7656 11169 7665 11203
rect 7665 11169 7699 11203
rect 7699 11169 7708 11203
rect 7656 11160 7708 11169
rect 7840 11160 7892 11212
rect 7748 11092 7800 11144
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 5632 11067 5684 11076
rect 5632 11033 5641 11067
rect 5641 11033 5675 11067
rect 5675 11033 5684 11067
rect 5632 11024 5684 11033
rect 8576 11024 8628 11076
rect 11428 11160 11480 11212
rect 11888 11296 11940 11348
rect 15292 11296 15344 11348
rect 15660 11296 15712 11348
rect 18512 11296 18564 11348
rect 12348 11228 12400 11280
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 13268 11160 13320 11212
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 15936 11203 15988 11212
rect 15936 11169 15945 11203
rect 15945 11169 15979 11203
rect 15979 11169 15988 11203
rect 15936 11160 15988 11169
rect 16304 11160 16356 11212
rect 18328 11160 18380 11212
rect 19248 11160 19300 11212
rect 22652 11160 22704 11212
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 16396 11092 16448 11144
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 21548 11092 21600 11144
rect 23296 11092 23348 11144
rect 23388 11092 23440 11144
rect 12624 11024 12676 11076
rect 16488 11067 16540 11076
rect 16488 11033 16497 11067
rect 16497 11033 16531 11067
rect 16531 11033 16540 11067
rect 16488 11024 16540 11033
rect 21364 11024 21416 11076
rect 21456 11067 21508 11076
rect 21456 11033 21465 11067
rect 21465 11033 21499 11067
rect 21499 11033 21508 11067
rect 21456 11024 21508 11033
rect 17684 10956 17736 11008
rect 18328 10999 18380 11008
rect 18328 10965 18337 10999
rect 18337 10965 18371 10999
rect 18371 10965 18380 10999
rect 18328 10956 18380 10965
rect 23020 10956 23072 11008
rect 4473 10854 4525 10906
rect 4537 10854 4589 10906
rect 4601 10854 4653 10906
rect 4665 10854 4717 10906
rect 4729 10854 4781 10906
rect 10200 10854 10252 10906
rect 10264 10854 10316 10906
rect 10328 10854 10380 10906
rect 10392 10854 10444 10906
rect 10456 10854 10508 10906
rect 15927 10854 15979 10906
rect 15991 10854 16043 10906
rect 16055 10854 16107 10906
rect 16119 10854 16171 10906
rect 16183 10854 16235 10906
rect 21654 10854 21706 10906
rect 21718 10854 21770 10906
rect 21782 10854 21834 10906
rect 21846 10854 21898 10906
rect 21910 10854 21962 10906
rect 5632 10752 5684 10804
rect 13728 10752 13780 10804
rect 13544 10684 13596 10736
rect 4804 10616 4856 10668
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 5080 10591 5132 10600
rect 5080 10557 5089 10591
rect 5089 10557 5123 10591
rect 5123 10557 5132 10591
rect 5080 10548 5132 10557
rect 13544 10591 13596 10600
rect 13544 10557 13553 10591
rect 13553 10557 13587 10591
rect 13587 10557 13596 10591
rect 13544 10548 13596 10557
rect 5448 10523 5500 10532
rect 5448 10489 5457 10523
rect 5457 10489 5491 10523
rect 5491 10489 5500 10523
rect 5448 10480 5500 10489
rect 18328 10752 18380 10804
rect 18420 10795 18472 10804
rect 18420 10761 18429 10795
rect 18429 10761 18463 10795
rect 18463 10761 18472 10795
rect 18420 10752 18472 10761
rect 18696 10752 18748 10804
rect 15292 10727 15344 10736
rect 15292 10693 15301 10727
rect 15301 10693 15335 10727
rect 15335 10693 15344 10727
rect 15292 10684 15344 10693
rect 15752 10684 15804 10736
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 21640 10616 21692 10668
rect 22100 10616 22152 10668
rect 19156 10548 19208 10600
rect 20904 10548 20956 10600
rect 21548 10591 21600 10600
rect 21548 10557 21557 10591
rect 21557 10557 21591 10591
rect 21591 10557 21600 10591
rect 21548 10548 21600 10557
rect 22008 10548 22060 10600
rect 23204 10591 23256 10600
rect 23204 10557 23213 10591
rect 23213 10557 23247 10591
rect 23247 10557 23256 10591
rect 23204 10548 23256 10557
rect 15936 10480 15988 10532
rect 19616 10480 19668 10532
rect 848 10412 900 10464
rect 5264 10412 5316 10464
rect 14280 10455 14332 10464
rect 14280 10421 14289 10455
rect 14289 10421 14323 10455
rect 14323 10421 14332 10455
rect 14280 10412 14332 10421
rect 15844 10412 15896 10464
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 19984 10455 20036 10464
rect 19984 10421 19993 10455
rect 19993 10421 20027 10455
rect 20027 10421 20036 10455
rect 19984 10412 20036 10421
rect 20444 10412 20496 10464
rect 22652 10455 22704 10464
rect 22652 10421 22661 10455
rect 22661 10421 22695 10455
rect 22695 10421 22704 10455
rect 22652 10412 22704 10421
rect 3813 10310 3865 10362
rect 3877 10310 3929 10362
rect 3941 10310 3993 10362
rect 4005 10310 4057 10362
rect 4069 10310 4121 10362
rect 9540 10310 9592 10362
rect 9604 10310 9656 10362
rect 9668 10310 9720 10362
rect 9732 10310 9784 10362
rect 9796 10310 9848 10362
rect 15267 10310 15319 10362
rect 15331 10310 15383 10362
rect 15395 10310 15447 10362
rect 15459 10310 15511 10362
rect 15523 10310 15575 10362
rect 20994 10310 21046 10362
rect 21058 10310 21110 10362
rect 21122 10310 21174 10362
rect 21186 10310 21238 10362
rect 21250 10310 21302 10362
rect 13544 10208 13596 10260
rect 18144 10208 18196 10260
rect 20904 10208 20956 10260
rect 21456 10208 21508 10260
rect 22008 10251 22060 10260
rect 22008 10217 22017 10251
rect 22017 10217 22051 10251
rect 22051 10217 22060 10251
rect 22008 10208 22060 10217
rect 22100 10251 22152 10260
rect 22100 10217 22109 10251
rect 22109 10217 22143 10251
rect 22143 10217 22152 10251
rect 22100 10208 22152 10217
rect 5080 10072 5132 10124
rect 8576 10140 8628 10192
rect 14280 10140 14332 10192
rect 20260 10140 20312 10192
rect 8208 10072 8260 10124
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 16396 10072 16448 10124
rect 18512 10072 18564 10124
rect 19248 10072 19300 10124
rect 19984 10072 20036 10124
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 7380 10004 7432 10056
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 16120 10004 16172 10056
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 19616 10047 19668 10056
rect 19616 10013 19625 10047
rect 19625 10013 19659 10047
rect 19659 10013 19668 10047
rect 19616 10004 19668 10013
rect 20444 10047 20496 10056
rect 20444 10013 20453 10047
rect 20453 10013 20487 10047
rect 20487 10013 20496 10047
rect 20444 10004 20496 10013
rect 1400 9911 1452 9920
rect 1400 9877 1409 9911
rect 1409 9877 1443 9911
rect 1443 9877 1452 9911
rect 1400 9868 1452 9877
rect 4896 9911 4948 9920
rect 4896 9877 4905 9911
rect 4905 9877 4939 9911
rect 4939 9877 4948 9911
rect 4896 9868 4948 9877
rect 7288 9868 7340 9920
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 19340 9936 19392 9988
rect 20720 10072 20772 10124
rect 22192 10140 22244 10192
rect 22652 10072 22704 10124
rect 23020 10115 23072 10124
rect 23020 10081 23029 10115
rect 23029 10081 23063 10115
rect 23063 10081 23072 10115
rect 23020 10072 23072 10081
rect 23112 10115 23164 10124
rect 23112 10081 23121 10115
rect 23121 10081 23155 10115
rect 23155 10081 23164 10115
rect 23112 10072 23164 10081
rect 21640 10047 21692 10056
rect 21640 10013 21649 10047
rect 21649 10013 21683 10047
rect 21683 10013 21692 10047
rect 21640 10004 21692 10013
rect 21548 9936 21600 9988
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 17868 9911 17920 9920
rect 17868 9877 17877 9911
rect 17877 9877 17911 9911
rect 17911 9877 17920 9911
rect 17868 9868 17920 9877
rect 17960 9868 18012 9920
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 23296 9868 23348 9920
rect 4473 9766 4525 9818
rect 4537 9766 4589 9818
rect 4601 9766 4653 9818
rect 4665 9766 4717 9818
rect 4729 9766 4781 9818
rect 10200 9766 10252 9818
rect 10264 9766 10316 9818
rect 10328 9766 10380 9818
rect 10392 9766 10444 9818
rect 10456 9766 10508 9818
rect 15927 9766 15979 9818
rect 15991 9766 16043 9818
rect 16055 9766 16107 9818
rect 16119 9766 16171 9818
rect 16183 9766 16235 9818
rect 21654 9766 21706 9818
rect 21718 9766 21770 9818
rect 21782 9766 21834 9818
rect 21846 9766 21898 9818
rect 21910 9766 21962 9818
rect 4896 9707 4948 9716
rect 4896 9673 4905 9707
rect 4905 9673 4939 9707
rect 4939 9673 4948 9707
rect 4896 9664 4948 9673
rect 7288 9664 7340 9716
rect 15384 9664 15436 9716
rect 4988 9639 5040 9648
rect 4988 9605 4997 9639
rect 4997 9605 5031 9639
rect 5031 9605 5040 9639
rect 4988 9596 5040 9605
rect 7380 9596 7432 9648
rect 13728 9596 13780 9648
rect 13820 9596 13872 9648
rect 17868 9664 17920 9716
rect 23572 9664 23624 9716
rect 17684 9596 17736 9648
rect 4988 9460 5040 9512
rect 8024 9460 8076 9512
rect 10600 9528 10652 9580
rect 10784 9528 10836 9580
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 10692 9460 10744 9512
rect 10876 9460 10928 9512
rect 11244 9392 11296 9444
rect 13360 9503 13412 9512
rect 13360 9469 13369 9503
rect 13369 9469 13403 9503
rect 13403 9469 13412 9503
rect 13360 9460 13412 9469
rect 16580 9528 16632 9580
rect 17960 9571 18012 9580
rect 15752 9460 15804 9512
rect 17960 9537 17969 9571
rect 17969 9537 18003 9571
rect 18003 9537 18012 9571
rect 17960 9528 18012 9537
rect 23664 9435 23716 9444
rect 23664 9401 23673 9435
rect 23673 9401 23707 9435
rect 23707 9401 23716 9435
rect 23664 9392 23716 9401
rect 4804 9324 4856 9376
rect 7380 9324 7432 9376
rect 9404 9324 9456 9376
rect 10876 9324 10928 9376
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 15660 9324 15712 9376
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16212 9324 16264 9333
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 3813 9222 3865 9274
rect 3877 9222 3929 9274
rect 3941 9222 3993 9274
rect 4005 9222 4057 9274
rect 4069 9222 4121 9274
rect 9540 9222 9592 9274
rect 9604 9222 9656 9274
rect 9668 9222 9720 9274
rect 9732 9222 9784 9274
rect 9796 9222 9848 9274
rect 15267 9222 15319 9274
rect 15331 9222 15383 9274
rect 15395 9222 15447 9274
rect 15459 9222 15511 9274
rect 15523 9222 15575 9274
rect 20994 9222 21046 9274
rect 21058 9222 21110 9274
rect 21122 9222 21174 9274
rect 21186 9222 21238 9274
rect 21250 9222 21302 9274
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 8576 9120 8628 9172
rect 10968 9120 11020 9172
rect 13360 9120 13412 9172
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 848 9052 900 9104
rect 8576 9027 8628 9036
rect 8576 8993 8585 9027
rect 8585 8993 8619 9027
rect 8619 8993 8628 9027
rect 8576 8984 8628 8993
rect 12808 9052 12860 9104
rect 14648 9052 14700 9104
rect 9404 8916 9456 8968
rect 10600 8848 10652 8900
rect 10968 8848 11020 8900
rect 11152 8916 11204 8968
rect 13912 8984 13964 9036
rect 16212 9027 16264 9036
rect 16212 8993 16221 9027
rect 16221 8993 16255 9027
rect 16255 8993 16264 9027
rect 16212 8984 16264 8993
rect 16396 9027 16448 9036
rect 16396 8993 16405 9027
rect 16405 8993 16439 9027
rect 16439 8993 16448 9027
rect 16396 8984 16448 8993
rect 19248 8984 19300 9036
rect 13728 8916 13780 8968
rect 17408 8916 17460 8968
rect 16304 8848 16356 8900
rect 10692 8780 10744 8832
rect 11980 8823 12032 8832
rect 11980 8789 11989 8823
rect 11989 8789 12023 8823
rect 12023 8789 12032 8823
rect 11980 8780 12032 8789
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 23664 8823 23716 8832
rect 23664 8789 23673 8823
rect 23673 8789 23707 8823
rect 23707 8789 23716 8823
rect 23664 8780 23716 8789
rect 4473 8678 4525 8730
rect 4537 8678 4589 8730
rect 4601 8678 4653 8730
rect 4665 8678 4717 8730
rect 4729 8678 4781 8730
rect 10200 8678 10252 8730
rect 10264 8678 10316 8730
rect 10328 8678 10380 8730
rect 10392 8678 10444 8730
rect 10456 8678 10508 8730
rect 15927 8678 15979 8730
rect 15991 8678 16043 8730
rect 16055 8678 16107 8730
rect 16119 8678 16171 8730
rect 16183 8678 16235 8730
rect 21654 8678 21706 8730
rect 21718 8678 21770 8730
rect 21782 8678 21834 8730
rect 21846 8678 21898 8730
rect 21910 8678 21962 8730
rect 5448 8576 5500 8628
rect 10876 8576 10928 8628
rect 13452 8576 13504 8628
rect 17408 8576 17460 8628
rect 16856 8508 16908 8560
rect 5632 8440 5684 8492
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 10784 8440 10836 8492
rect 11244 8440 11296 8492
rect 13912 8440 13964 8492
rect 15660 8440 15712 8492
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 4344 8347 4396 8356
rect 4344 8313 4353 8347
rect 4353 8313 4387 8347
rect 4387 8313 4396 8347
rect 4344 8304 4396 8313
rect 10600 8304 10652 8356
rect 11152 8372 11204 8424
rect 11980 8372 12032 8424
rect 13636 8415 13688 8424
rect 13636 8381 13645 8415
rect 13645 8381 13679 8415
rect 13679 8381 13688 8415
rect 13636 8372 13688 8381
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 16396 8372 16448 8424
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 19248 8415 19300 8424
rect 19248 8381 19257 8415
rect 19257 8381 19291 8415
rect 19291 8381 19300 8415
rect 19248 8372 19300 8381
rect 22560 8440 22612 8492
rect 22468 8415 22520 8424
rect 22468 8381 22477 8415
rect 22477 8381 22511 8415
rect 22511 8381 22520 8415
rect 22468 8372 22520 8381
rect 22928 8483 22980 8492
rect 22928 8449 22962 8483
rect 22962 8449 22980 8483
rect 22928 8440 22980 8449
rect 12348 8304 12400 8356
rect 17960 8304 18012 8356
rect 4252 8236 4304 8288
rect 5172 8236 5224 8288
rect 10508 8236 10560 8288
rect 20720 8304 20772 8356
rect 23388 8304 23440 8356
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 21732 8236 21784 8288
rect 22192 8236 22244 8288
rect 23020 8236 23072 8288
rect 3813 8134 3865 8186
rect 3877 8134 3929 8186
rect 3941 8134 3993 8186
rect 4005 8134 4057 8186
rect 4069 8134 4121 8186
rect 9540 8134 9592 8186
rect 9604 8134 9656 8186
rect 9668 8134 9720 8186
rect 9732 8134 9784 8186
rect 9796 8134 9848 8186
rect 15267 8134 15319 8186
rect 15331 8134 15383 8186
rect 15395 8134 15447 8186
rect 15459 8134 15511 8186
rect 15523 8134 15575 8186
rect 20994 8134 21046 8186
rect 21058 8134 21110 8186
rect 21122 8134 21174 8186
rect 21186 8134 21238 8186
rect 21250 8134 21302 8186
rect 5632 8075 5684 8084
rect 5632 8041 5641 8075
rect 5641 8041 5675 8075
rect 5675 8041 5684 8075
rect 5632 8032 5684 8041
rect 10232 8032 10284 8084
rect 13636 8032 13688 8084
rect 13912 8075 13964 8084
rect 13912 8041 13921 8075
rect 13921 8041 13955 8075
rect 13955 8041 13964 8075
rect 13912 8032 13964 8041
rect 15844 8032 15896 8084
rect 16672 8032 16724 8084
rect 22100 8032 22152 8084
rect 22468 8032 22520 8084
rect 10048 7964 10100 8016
rect 15660 7964 15712 8016
rect 4528 7896 4580 7948
rect 848 7828 900 7880
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 4896 7896 4948 7948
rect 5080 7896 5132 7948
rect 5356 7896 5408 7948
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 11152 7896 11204 7948
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 13544 7939 13596 7948
rect 5724 7828 5776 7880
rect 7288 7828 7340 7880
rect 10692 7828 10744 7880
rect 13544 7905 13553 7939
rect 13553 7905 13587 7939
rect 13587 7905 13596 7939
rect 13544 7896 13596 7905
rect 14648 7939 14700 7948
rect 14648 7905 14657 7939
rect 14657 7905 14691 7939
rect 14691 7905 14700 7939
rect 14648 7896 14700 7905
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 21364 7964 21416 8016
rect 16580 7896 16632 7948
rect 16948 7896 17000 7948
rect 20904 7939 20956 7948
rect 20904 7905 20913 7939
rect 20913 7905 20947 7939
rect 20947 7905 20956 7939
rect 20904 7896 20956 7905
rect 2596 7692 2648 7744
rect 5080 7735 5132 7744
rect 5080 7701 5089 7735
rect 5089 7701 5123 7735
rect 5123 7701 5132 7735
rect 5080 7692 5132 7701
rect 5172 7735 5224 7744
rect 5172 7701 5181 7735
rect 5181 7701 5215 7735
rect 5215 7701 5224 7735
rect 5172 7692 5224 7701
rect 7104 7760 7156 7812
rect 13176 7760 13228 7812
rect 16672 7828 16724 7880
rect 21732 7939 21784 7948
rect 21732 7905 21741 7939
rect 21741 7905 21775 7939
rect 21775 7905 21784 7939
rect 21732 7896 21784 7905
rect 14464 7803 14516 7812
rect 14464 7769 14473 7803
rect 14473 7769 14507 7803
rect 14507 7769 14516 7803
rect 14464 7760 14516 7769
rect 14556 7735 14608 7744
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 15200 7760 15252 7812
rect 16488 7692 16540 7744
rect 21088 7692 21140 7744
rect 21548 7760 21600 7812
rect 23112 7939 23164 7948
rect 23112 7905 23121 7939
rect 23121 7905 23155 7939
rect 23155 7905 23164 7939
rect 23112 7896 23164 7905
rect 22192 7828 22244 7880
rect 23480 7871 23532 7880
rect 22008 7760 22060 7812
rect 23480 7837 23514 7871
rect 23514 7837 23532 7871
rect 23480 7828 23532 7837
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 4473 7590 4525 7642
rect 4537 7590 4589 7642
rect 4601 7590 4653 7642
rect 4665 7590 4717 7642
rect 4729 7590 4781 7642
rect 10200 7590 10252 7642
rect 10264 7590 10316 7642
rect 10328 7590 10380 7642
rect 10392 7590 10444 7642
rect 10456 7590 10508 7642
rect 15927 7590 15979 7642
rect 15991 7590 16043 7642
rect 16055 7590 16107 7642
rect 16119 7590 16171 7642
rect 16183 7590 16235 7642
rect 21654 7590 21706 7642
rect 21718 7590 21770 7642
rect 21782 7590 21834 7642
rect 21846 7590 21898 7642
rect 21910 7590 21962 7642
rect 2596 7420 2648 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 4344 7488 4396 7540
rect 5080 7488 5132 7540
rect 7288 7531 7340 7540
rect 7288 7497 7297 7531
rect 7297 7497 7331 7531
rect 7331 7497 7340 7531
rect 7288 7488 7340 7497
rect 13268 7488 13320 7540
rect 14556 7488 14608 7540
rect 22560 7531 22612 7540
rect 22560 7497 22569 7531
rect 22569 7497 22603 7531
rect 22603 7497 22612 7531
rect 22560 7488 22612 7497
rect 22928 7531 22980 7540
rect 22928 7497 22937 7531
rect 22937 7497 22971 7531
rect 22971 7497 22980 7531
rect 22928 7488 22980 7497
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 4252 7327 4304 7336
rect 4252 7293 4261 7327
rect 4261 7293 4295 7327
rect 4295 7293 4304 7327
rect 4252 7284 4304 7293
rect 4804 7216 4856 7268
rect 5356 7352 5408 7404
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 7472 7352 7524 7404
rect 5264 7216 5316 7268
rect 7932 7284 7984 7336
rect 8208 7284 8260 7336
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 9312 7352 9364 7404
rect 14464 7352 14516 7404
rect 15200 7352 15252 7404
rect 15568 7352 15620 7404
rect 16304 7352 16356 7404
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 21364 7352 21416 7404
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 23664 7352 23716 7361
rect 18880 7284 18932 7336
rect 19064 7327 19116 7336
rect 19064 7293 19073 7327
rect 19073 7293 19107 7327
rect 19107 7293 19116 7327
rect 19064 7284 19116 7293
rect 21088 7327 21140 7336
rect 21088 7293 21097 7327
rect 21097 7293 21131 7327
rect 21131 7293 21140 7327
rect 21088 7284 21140 7293
rect 22008 7284 22060 7336
rect 22100 7327 22152 7336
rect 22100 7293 22109 7327
rect 22109 7293 22143 7327
rect 22143 7293 22152 7327
rect 22100 7284 22152 7293
rect 23204 7327 23256 7336
rect 23204 7293 23213 7327
rect 23213 7293 23247 7327
rect 23247 7293 23256 7327
rect 23204 7284 23256 7293
rect 16396 7216 16448 7268
rect 5448 7148 5500 7200
rect 7012 7148 7064 7200
rect 8024 7191 8076 7200
rect 8024 7157 8033 7191
rect 8033 7157 8067 7191
rect 8067 7157 8076 7191
rect 8024 7148 8076 7157
rect 8392 7148 8444 7200
rect 9312 7148 9364 7200
rect 17040 7148 17092 7200
rect 3813 7046 3865 7098
rect 3877 7046 3929 7098
rect 3941 7046 3993 7098
rect 4005 7046 4057 7098
rect 4069 7046 4121 7098
rect 9540 7046 9592 7098
rect 9604 7046 9656 7098
rect 9668 7046 9720 7098
rect 9732 7046 9784 7098
rect 9796 7046 9848 7098
rect 15267 7046 15319 7098
rect 15331 7046 15383 7098
rect 15395 7046 15447 7098
rect 15459 7046 15511 7098
rect 15523 7046 15575 7098
rect 20994 7046 21046 7098
rect 21058 7046 21110 7098
rect 21122 7046 21174 7098
rect 21186 7046 21238 7098
rect 21250 7046 21302 7098
rect 5172 6944 5224 6996
rect 5264 6944 5316 6996
rect 5448 6944 5500 6996
rect 7472 6987 7524 6996
rect 7472 6953 7481 6987
rect 7481 6953 7515 6987
rect 7515 6953 7524 6987
rect 7472 6944 7524 6953
rect 16304 6987 16356 6996
rect 16304 6953 16313 6987
rect 16313 6953 16347 6987
rect 16347 6953 16356 6987
rect 16304 6944 16356 6953
rect 4344 6876 4396 6928
rect 4804 6808 4856 6860
rect 4988 6808 5040 6860
rect 8576 6808 8628 6860
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 7380 6740 7432 6792
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8760 6740 8812 6792
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 10968 6740 11020 6792
rect 13544 6876 13596 6928
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 18144 6876 18196 6928
rect 19248 6876 19300 6928
rect 21548 6876 21600 6928
rect 22192 6919 22244 6928
rect 22192 6885 22201 6919
rect 22201 6885 22235 6919
rect 22235 6885 22244 6919
rect 22192 6876 22244 6885
rect 18696 6808 18748 6860
rect 22100 6808 22152 6860
rect 13176 6740 13228 6792
rect 18880 6783 18932 6792
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 18880 6740 18932 6749
rect 22468 6740 22520 6792
rect 23572 6740 23624 6792
rect 15660 6672 15712 6724
rect 7012 6604 7064 6656
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 9956 6604 10008 6656
rect 13452 6604 13504 6656
rect 15200 6604 15252 6656
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 16672 6647 16724 6656
rect 16672 6613 16681 6647
rect 16681 6613 16715 6647
rect 16715 6613 16724 6647
rect 16672 6604 16724 6613
rect 17224 6604 17276 6656
rect 18512 6604 18564 6656
rect 23664 6647 23716 6656
rect 23664 6613 23673 6647
rect 23673 6613 23707 6647
rect 23707 6613 23716 6647
rect 23664 6604 23716 6613
rect 4473 6502 4525 6554
rect 4537 6502 4589 6554
rect 4601 6502 4653 6554
rect 4665 6502 4717 6554
rect 4729 6502 4781 6554
rect 10200 6502 10252 6554
rect 10264 6502 10316 6554
rect 10328 6502 10380 6554
rect 10392 6502 10444 6554
rect 10456 6502 10508 6554
rect 15927 6502 15979 6554
rect 15991 6502 16043 6554
rect 16055 6502 16107 6554
rect 16119 6502 16171 6554
rect 16183 6502 16235 6554
rect 21654 6502 21706 6554
rect 21718 6502 21770 6554
rect 21782 6502 21834 6554
rect 21846 6502 21898 6554
rect 21910 6502 21962 6554
rect 9588 6400 9640 6452
rect 10692 6400 10744 6452
rect 10876 6400 10928 6452
rect 10968 6443 11020 6452
rect 10968 6409 10977 6443
rect 10977 6409 11011 6443
rect 11011 6409 11020 6443
rect 10968 6400 11020 6409
rect 13544 6400 13596 6452
rect 15476 6400 15528 6452
rect 18236 6400 18288 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 8760 6332 8812 6384
rect 8484 6264 8536 6316
rect 4988 6196 5040 6248
rect 8300 6196 8352 6248
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 8668 6196 8720 6248
rect 14280 6332 14332 6384
rect 18512 6375 18564 6384
rect 18512 6341 18521 6375
rect 18521 6341 18555 6375
rect 18555 6341 18564 6375
rect 18512 6332 18564 6341
rect 19248 6332 19300 6384
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 8392 6128 8444 6180
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 12716 6239 12768 6248
rect 12716 6205 12725 6239
rect 12725 6205 12759 6239
rect 12759 6205 12768 6239
rect 12716 6196 12768 6205
rect 13268 6196 13320 6248
rect 13820 6264 13872 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 18972 6264 19024 6316
rect 19156 6307 19208 6316
rect 19156 6273 19165 6307
rect 19165 6273 19199 6307
rect 19199 6273 19208 6307
rect 19156 6264 19208 6273
rect 14372 6196 14424 6248
rect 18144 6196 18196 6248
rect 19248 6239 19300 6248
rect 19248 6205 19257 6239
rect 19257 6205 19291 6239
rect 19291 6205 19300 6239
rect 19248 6196 19300 6205
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 19984 6264 20036 6273
rect 23664 6307 23716 6316
rect 23664 6273 23673 6307
rect 23673 6273 23707 6307
rect 23707 6273 23716 6307
rect 23664 6264 23716 6273
rect 20168 6196 20220 6248
rect 7932 6060 7984 6112
rect 18880 6128 18932 6180
rect 13360 6060 13412 6112
rect 15844 6060 15896 6112
rect 17592 6060 17644 6112
rect 3813 5958 3865 6010
rect 3877 5958 3929 6010
rect 3941 5958 3993 6010
rect 4005 5958 4057 6010
rect 4069 5958 4121 6010
rect 9540 5958 9592 6010
rect 9604 5958 9656 6010
rect 9668 5958 9720 6010
rect 9732 5958 9784 6010
rect 9796 5958 9848 6010
rect 15267 5958 15319 6010
rect 15331 5958 15383 6010
rect 15395 5958 15447 6010
rect 15459 5958 15511 6010
rect 15523 5958 15575 6010
rect 20994 5958 21046 6010
rect 21058 5958 21110 6010
rect 21122 5958 21174 6010
rect 21186 5958 21238 6010
rect 21250 5958 21302 6010
rect 7380 5856 7432 5908
rect 8668 5899 8720 5908
rect 8668 5865 8677 5899
rect 8677 5865 8711 5899
rect 8711 5865 8720 5899
rect 8668 5856 8720 5865
rect 10876 5856 10928 5908
rect 12716 5856 12768 5908
rect 17224 5899 17276 5908
rect 17224 5865 17233 5899
rect 17233 5865 17267 5899
rect 17267 5865 17276 5899
rect 17224 5856 17276 5865
rect 19156 5856 19208 5908
rect 19248 5856 19300 5908
rect 23296 5856 23348 5908
rect 4988 5763 5040 5772
rect 4988 5729 4997 5763
rect 4997 5729 5031 5763
rect 5031 5729 5040 5763
rect 4988 5720 5040 5729
rect 5540 5652 5592 5704
rect 10600 5652 10652 5704
rect 10876 5720 10928 5772
rect 14280 5788 14332 5840
rect 18972 5788 19024 5840
rect 13268 5720 13320 5772
rect 14372 5720 14424 5772
rect 18052 5720 18104 5772
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 19984 5652 20036 5704
rect 23388 5652 23440 5704
rect 20168 5584 20220 5636
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 11520 5516 11572 5525
rect 13820 5516 13872 5568
rect 4473 5414 4525 5466
rect 4537 5414 4589 5466
rect 4601 5414 4653 5466
rect 4665 5414 4717 5466
rect 4729 5414 4781 5466
rect 10200 5414 10252 5466
rect 10264 5414 10316 5466
rect 10328 5414 10380 5466
rect 10392 5414 10444 5466
rect 10456 5414 10508 5466
rect 15927 5414 15979 5466
rect 15991 5414 16043 5466
rect 16055 5414 16107 5466
rect 16119 5414 16171 5466
rect 16183 5414 16235 5466
rect 21654 5414 21706 5466
rect 21718 5414 21770 5466
rect 21782 5414 21834 5466
rect 21846 5414 21898 5466
rect 21910 5414 21962 5466
rect 5080 5355 5132 5364
rect 5080 5321 5089 5355
rect 5089 5321 5123 5355
rect 5123 5321 5132 5355
rect 5080 5312 5132 5321
rect 5540 5355 5592 5364
rect 5540 5321 5549 5355
rect 5549 5321 5583 5355
rect 5583 5321 5592 5355
rect 5540 5312 5592 5321
rect 14372 5355 14424 5364
rect 14372 5321 14381 5355
rect 14381 5321 14415 5355
rect 14415 5321 14424 5355
rect 14372 5312 14424 5321
rect 14924 5312 14976 5364
rect 5356 5244 5408 5296
rect 4344 5176 4396 5228
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 4896 5108 4948 5160
rect 7656 5108 7708 5160
rect 8300 5108 8352 5160
rect 11520 5244 11572 5296
rect 11336 5176 11388 5228
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 14832 5108 14884 5160
rect 17868 5219 17920 5228
rect 17868 5185 17877 5219
rect 17877 5185 17911 5219
rect 17911 5185 17920 5219
rect 17868 5176 17920 5185
rect 15752 5151 15804 5160
rect 15752 5117 15761 5151
rect 15761 5117 15795 5151
rect 15795 5117 15804 5151
rect 15752 5108 15804 5117
rect 17500 5108 17552 5160
rect 18052 5108 18104 5160
rect 19984 5312 20036 5364
rect 20168 5312 20220 5364
rect 20812 5176 20864 5228
rect 21364 5176 21416 5228
rect 23664 5219 23716 5228
rect 23664 5185 23673 5219
rect 23673 5185 23707 5219
rect 23707 5185 23716 5219
rect 23664 5176 23716 5185
rect 20352 5151 20404 5160
rect 20352 5117 20361 5151
rect 20361 5117 20395 5151
rect 20395 5117 20404 5151
rect 20352 5108 20404 5117
rect 20444 5151 20496 5160
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 20904 5108 20956 5160
rect 21456 5108 21508 5160
rect 23112 5108 23164 5160
rect 8576 5015 8628 5024
rect 8576 4981 8585 5015
rect 8585 4981 8619 5015
rect 8619 4981 8628 5015
rect 8576 4972 8628 4981
rect 15752 4972 15804 5024
rect 3813 4870 3865 4922
rect 3877 4870 3929 4922
rect 3941 4870 3993 4922
rect 4005 4870 4057 4922
rect 4069 4870 4121 4922
rect 9540 4870 9592 4922
rect 9604 4870 9656 4922
rect 9668 4870 9720 4922
rect 9732 4870 9784 4922
rect 9796 4870 9848 4922
rect 15267 4870 15319 4922
rect 15331 4870 15383 4922
rect 15395 4870 15447 4922
rect 15459 4870 15511 4922
rect 15523 4870 15575 4922
rect 20994 4870 21046 4922
rect 21058 4870 21110 4922
rect 21122 4870 21174 4922
rect 21186 4870 21238 4922
rect 21250 4870 21302 4922
rect 5448 4768 5500 4820
rect 10876 4811 10928 4820
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 14556 4768 14608 4820
rect 20352 4768 20404 4820
rect 20904 4768 20956 4820
rect 7288 4700 7340 4752
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 5632 4564 5684 4616
rect 8576 4632 8628 4684
rect 15752 4700 15804 4752
rect 21548 4632 21600 4684
rect 4160 4496 4212 4548
rect 7472 4539 7524 4548
rect 7472 4505 7481 4539
rect 7481 4505 7515 4539
rect 7515 4505 7524 4539
rect 7472 4496 7524 4505
rect 7564 4496 7616 4548
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 14832 4564 14884 4616
rect 10600 4496 10652 4548
rect 21364 4564 21416 4616
rect 23480 4564 23532 4616
rect 23664 4607 23716 4616
rect 23664 4573 23673 4607
rect 23673 4573 23707 4607
rect 23707 4573 23716 4607
rect 23664 4564 23716 4573
rect 20904 4496 20956 4548
rect 4988 4471 5040 4480
rect 4988 4437 4997 4471
rect 4997 4437 5031 4471
rect 5031 4437 5040 4471
rect 4988 4428 5040 4437
rect 5172 4428 5224 4480
rect 8116 4428 8168 4480
rect 4473 4326 4525 4378
rect 4537 4326 4589 4378
rect 4601 4326 4653 4378
rect 4665 4326 4717 4378
rect 4729 4326 4781 4378
rect 10200 4326 10252 4378
rect 10264 4326 10316 4378
rect 10328 4326 10380 4378
rect 10392 4326 10444 4378
rect 10456 4326 10508 4378
rect 15927 4326 15979 4378
rect 15991 4326 16043 4378
rect 16055 4326 16107 4378
rect 16119 4326 16171 4378
rect 16183 4326 16235 4378
rect 21654 4326 21706 4378
rect 21718 4326 21770 4378
rect 21782 4326 21834 4378
rect 21846 4326 21898 4378
rect 21910 4326 21962 4378
rect 4344 4224 4396 4276
rect 4804 4224 4856 4276
rect 7472 4224 7524 4276
rect 8116 4267 8168 4276
rect 8116 4233 8125 4267
rect 8125 4233 8159 4267
rect 8159 4233 8168 4267
rect 8116 4224 8168 4233
rect 11152 4224 11204 4276
rect 18144 4224 18196 4276
rect 10600 4156 10652 4208
rect 4160 4088 4212 4140
rect 4896 4088 4948 4140
rect 5816 4088 5868 4140
rect 7288 4131 7340 4140
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 10692 4131 10744 4140
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 7564 4020 7616 4072
rect 7656 4063 7708 4072
rect 7656 4029 7665 4063
rect 7665 4029 7699 4063
rect 7699 4029 7708 4063
rect 7656 4020 7708 4029
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 7932 4020 7984 4072
rect 4804 3952 4856 4004
rect 4896 3884 4948 3936
rect 8484 3995 8536 4004
rect 8484 3961 8493 3995
rect 8493 3961 8527 3995
rect 8527 3961 8536 3995
rect 8484 3952 8536 3961
rect 10048 3952 10100 4004
rect 14832 4020 14884 4072
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 15844 4063 15896 4072
rect 15844 4029 15853 4063
rect 15853 4029 15887 4063
rect 15887 4029 15896 4063
rect 15844 4020 15896 4029
rect 17592 4131 17644 4140
rect 17592 4097 17601 4131
rect 17601 4097 17635 4131
rect 17635 4097 17644 4131
rect 17592 4088 17644 4097
rect 15568 3995 15620 4004
rect 15568 3961 15577 3995
rect 15577 3961 15611 3995
rect 15611 3961 15620 3995
rect 15568 3952 15620 3961
rect 14832 3884 14884 3936
rect 16672 3952 16724 4004
rect 17684 4063 17736 4072
rect 17684 4029 17693 4063
rect 17693 4029 17727 4063
rect 17727 4029 17736 4063
rect 17684 4020 17736 4029
rect 18144 4088 18196 4140
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 18328 4063 18380 4072
rect 18328 4029 18337 4063
rect 18337 4029 18371 4063
rect 18371 4029 18380 4063
rect 18328 4020 18380 4029
rect 3813 3782 3865 3834
rect 3877 3782 3929 3834
rect 3941 3782 3993 3834
rect 4005 3782 4057 3834
rect 4069 3782 4121 3834
rect 9540 3782 9592 3834
rect 9604 3782 9656 3834
rect 9668 3782 9720 3834
rect 9732 3782 9784 3834
rect 9796 3782 9848 3834
rect 15267 3782 15319 3834
rect 15331 3782 15383 3834
rect 15395 3782 15447 3834
rect 15459 3782 15511 3834
rect 15523 3782 15575 3834
rect 20994 3782 21046 3834
rect 21058 3782 21110 3834
rect 21122 3782 21174 3834
rect 21186 3782 21238 3834
rect 21250 3782 21302 3834
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 7932 3723 7984 3732
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 10600 3723 10652 3732
rect 10600 3689 10609 3723
rect 10609 3689 10643 3723
rect 10643 3689 10652 3723
rect 10600 3680 10652 3689
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 14740 3723 14792 3732
rect 14740 3689 14749 3723
rect 14749 3689 14783 3723
rect 14783 3689 14792 3723
rect 14740 3680 14792 3689
rect 15200 3723 15252 3732
rect 15200 3689 15209 3723
rect 15209 3689 15243 3723
rect 15243 3689 15252 3723
rect 15200 3680 15252 3689
rect 17592 3680 17644 3732
rect 17684 3680 17736 3732
rect 18328 3723 18380 3732
rect 18328 3689 18337 3723
rect 18337 3689 18371 3723
rect 18371 3689 18380 3723
rect 18328 3680 18380 3689
rect 20904 3680 20956 3732
rect 4896 3476 4948 3528
rect 6920 3476 6972 3528
rect 7288 3476 7340 3528
rect 7656 3476 7708 3528
rect 11152 3544 11204 3596
rect 12532 3612 12584 3664
rect 13728 3612 13780 3664
rect 18144 3612 18196 3664
rect 12072 3587 12124 3596
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 12072 3544 12124 3553
rect 14832 3544 14884 3596
rect 17868 3544 17920 3596
rect 4804 3451 4856 3460
rect 4804 3417 4813 3451
rect 4813 3417 4847 3451
rect 4847 3417 4856 3451
rect 4804 3408 4856 3417
rect 9864 3408 9916 3460
rect 15844 3476 15896 3528
rect 21456 3544 21508 3596
rect 14832 3451 14884 3460
rect 14832 3417 14841 3451
rect 14841 3417 14875 3451
rect 14875 3417 14884 3451
rect 14832 3408 14884 3417
rect 18144 3451 18196 3460
rect 18144 3417 18153 3451
rect 18153 3417 18187 3451
rect 18187 3417 18196 3451
rect 18144 3408 18196 3417
rect 18236 3408 18288 3460
rect 23664 3519 23716 3528
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 19524 3408 19576 3460
rect 10048 3340 10100 3392
rect 11888 3383 11940 3392
rect 11888 3349 11897 3383
rect 11897 3349 11931 3383
rect 11931 3349 11940 3383
rect 11888 3340 11940 3349
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 4473 3238 4525 3290
rect 4537 3238 4589 3290
rect 4601 3238 4653 3290
rect 4665 3238 4717 3290
rect 4729 3238 4781 3290
rect 10200 3238 10252 3290
rect 10264 3238 10316 3290
rect 10328 3238 10380 3290
rect 10392 3238 10444 3290
rect 10456 3238 10508 3290
rect 15927 3238 15979 3290
rect 15991 3238 16043 3290
rect 16055 3238 16107 3290
rect 16119 3238 16171 3290
rect 16183 3238 16235 3290
rect 21654 3238 21706 3290
rect 21718 3238 21770 3290
rect 21782 3238 21834 3290
rect 21846 3238 21898 3290
rect 21910 3238 21962 3290
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 6920 3136 6972 3188
rect 7380 3136 7432 3188
rect 7656 3136 7708 3188
rect 10048 3136 10100 3188
rect 14832 3136 14884 3188
rect 15844 3136 15896 3188
rect 4160 3068 4212 3120
rect 4528 3043 4580 3052
rect 4528 3009 4572 3043
rect 4572 3009 4580 3043
rect 4528 3000 4580 3009
rect 6920 3000 6972 3052
rect 4252 2932 4304 2984
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 12072 3068 12124 3120
rect 16028 3068 16080 3120
rect 9864 3000 9916 3052
rect 14648 3000 14700 3052
rect 15016 3043 15068 3052
rect 15016 3009 15025 3043
rect 15025 3009 15059 3043
rect 15059 3009 15068 3043
rect 15016 3000 15068 3009
rect 15660 3000 15712 3052
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 13728 2864 13780 2916
rect 15936 2975 15988 2984
rect 15936 2941 15945 2975
rect 15945 2941 15979 2975
rect 15979 2941 15988 2975
rect 15936 2932 15988 2941
rect 18144 3136 18196 3188
rect 18788 3136 18840 3188
rect 23480 3179 23532 3188
rect 23480 3145 23489 3179
rect 23489 3145 23523 3179
rect 23523 3145 23532 3179
rect 23480 3136 23532 3145
rect 18236 2932 18288 2984
rect 19524 3000 19576 3052
rect 23664 3043 23716 3052
rect 23664 3009 23673 3043
rect 23673 3009 23707 3043
rect 23707 3009 23716 3043
rect 23664 3000 23716 3009
rect 19432 2932 19484 2984
rect 20444 2864 20496 2916
rect 4712 2796 4764 2848
rect 6828 2796 6880 2848
rect 15016 2796 15068 2848
rect 17500 2796 17552 2848
rect 3813 2694 3865 2746
rect 3877 2694 3929 2746
rect 3941 2694 3993 2746
rect 4005 2694 4057 2746
rect 4069 2694 4121 2746
rect 9540 2694 9592 2746
rect 9604 2694 9656 2746
rect 9668 2694 9720 2746
rect 9732 2694 9784 2746
rect 9796 2694 9848 2746
rect 15267 2694 15319 2746
rect 15331 2694 15383 2746
rect 15395 2694 15447 2746
rect 15459 2694 15511 2746
rect 15523 2694 15575 2746
rect 20994 2694 21046 2746
rect 21058 2694 21110 2746
rect 21122 2694 21174 2746
rect 21186 2694 21238 2746
rect 21250 2694 21302 2746
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 4528 2635 4580 2644
rect 4528 2601 4537 2635
rect 4537 2601 4571 2635
rect 4571 2601 4580 2635
rect 4528 2592 4580 2601
rect 4896 2592 4948 2644
rect 6920 2592 6972 2644
rect 7104 2592 7156 2644
rect 10968 2592 11020 2644
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 12624 2592 12676 2644
rect 13360 2592 13412 2644
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 15108 2592 15160 2644
rect 15936 2592 15988 2644
rect 16028 2592 16080 2644
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 19524 2592 19576 2644
rect 6828 2524 6880 2576
rect 7288 2567 7340 2576
rect 7288 2533 7297 2567
rect 7297 2533 7331 2567
rect 7331 2533 7340 2567
rect 7288 2524 7340 2533
rect 16488 2524 16540 2576
rect 17500 2567 17552 2576
rect 17500 2533 17509 2567
rect 17509 2533 17543 2567
rect 17543 2533 17552 2567
rect 17500 2524 17552 2533
rect 4712 2456 4764 2508
rect 5264 2499 5316 2508
rect 5264 2465 5273 2499
rect 5273 2465 5307 2499
rect 5307 2465 5316 2499
rect 5264 2456 5316 2465
rect 7196 2456 7248 2508
rect 3240 2388 3292 2440
rect 3884 2388 3936 2440
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 4528 2388 4580 2440
rect 5816 2388 5868 2440
rect 7012 2388 7064 2440
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 8024 2431 8076 2440
rect 8024 2397 8033 2431
rect 8033 2397 8067 2431
rect 8067 2397 8076 2431
rect 8024 2388 8076 2397
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10600 2388 10652 2440
rect 10968 2388 11020 2440
rect 11612 2388 11664 2440
rect 12256 2388 12308 2440
rect 12900 2388 12952 2440
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14188 2388 14240 2440
rect 15016 2431 15068 2440
rect 15016 2397 15050 2431
rect 15050 2397 15068 2431
rect 15016 2388 15068 2397
rect 15568 2388 15620 2440
rect 5172 2320 5224 2372
rect 10784 2320 10836 2372
rect 14832 2320 14884 2372
rect 15844 2388 15896 2440
rect 16396 2431 16448 2440
rect 16396 2397 16405 2431
rect 16405 2397 16439 2431
rect 16439 2397 16448 2431
rect 16396 2388 16448 2397
rect 17040 2431 17092 2440
rect 17040 2397 17049 2431
rect 17049 2397 17083 2431
rect 17083 2397 17092 2431
rect 17040 2388 17092 2397
rect 17408 2388 17460 2440
rect 17960 2388 18012 2440
rect 18696 2388 18748 2440
rect 19340 2388 19392 2440
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 20812 2388 20864 2440
rect 21272 2388 21324 2440
rect 6460 2252 6512 2304
rect 7748 2252 7800 2304
rect 8392 2252 8444 2304
rect 9036 2252 9088 2304
rect 9680 2252 9732 2304
rect 13544 2252 13596 2304
rect 15568 2252 15620 2304
rect 16304 2252 16356 2304
rect 16764 2252 16816 2304
rect 18052 2252 18104 2304
rect 19984 2252 20036 2304
rect 20628 2252 20680 2304
rect 4473 2150 4525 2202
rect 4537 2150 4589 2202
rect 4601 2150 4653 2202
rect 4665 2150 4717 2202
rect 4729 2150 4781 2202
rect 10200 2150 10252 2202
rect 10264 2150 10316 2202
rect 10328 2150 10380 2202
rect 10392 2150 10444 2202
rect 10456 2150 10508 2202
rect 15927 2150 15979 2202
rect 15991 2150 16043 2202
rect 16055 2150 16107 2202
rect 16119 2150 16171 2202
rect 16183 2150 16235 2202
rect 21654 2150 21706 2202
rect 21718 2150 21770 2202
rect 21782 2150 21834 2202
rect 21846 2150 21898 2202
rect 21910 2150 21962 2202
<< metal2 >>
rect 5814 26516 5870 27316
rect 6458 26516 6514 27316
rect 7102 26516 7158 27316
rect 7746 26516 7802 27316
rect 8390 26516 8446 27316
rect 9034 26516 9090 27316
rect 9678 26516 9734 27316
rect 10322 26516 10378 27316
rect 10428 26574 10640 26602
rect 4473 25052 4781 25061
rect 4473 25050 4479 25052
rect 4535 25050 4559 25052
rect 4615 25050 4639 25052
rect 4695 25050 4719 25052
rect 4775 25050 4781 25052
rect 4535 24998 4537 25050
rect 4717 24998 4719 25050
rect 4473 24996 4479 24998
rect 4535 24996 4559 24998
rect 4615 24996 4639 24998
rect 4695 24996 4719 24998
rect 4775 24996 4781 24998
rect 4473 24987 4781 24996
rect 5828 24818 5856 26516
rect 6472 24818 6500 26516
rect 7116 24818 7144 26516
rect 7760 24818 7788 26516
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 6460 24812 6512 24818
rect 6460 24754 6512 24760
rect 7104 24812 7156 24818
rect 7104 24754 7156 24760
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 8404 24682 8432 26516
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 6092 24608 6144 24614
rect 6092 24550 6144 24556
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 3813 24508 4121 24517
rect 3813 24506 3819 24508
rect 3875 24506 3899 24508
rect 3955 24506 3979 24508
rect 4035 24506 4059 24508
rect 4115 24506 4121 24508
rect 3875 24454 3877 24506
rect 4057 24454 4059 24506
rect 3813 24452 3819 24454
rect 3875 24452 3899 24454
rect 3955 24452 3979 24454
rect 4035 24452 4059 24454
rect 4115 24452 4121 24454
rect 3813 24443 4121 24452
rect 4473 23964 4781 23973
rect 4473 23962 4479 23964
rect 4535 23962 4559 23964
rect 4615 23962 4639 23964
rect 4695 23962 4719 23964
rect 4775 23962 4781 23964
rect 4535 23910 4537 23962
rect 4717 23910 4719 23962
rect 4473 23908 4479 23910
rect 4535 23908 4559 23910
rect 4615 23908 4639 23910
rect 4695 23908 4719 23910
rect 4775 23908 4781 23910
rect 4473 23899 4781 23908
rect 3813 23420 4121 23429
rect 3813 23418 3819 23420
rect 3875 23418 3899 23420
rect 3955 23418 3979 23420
rect 4035 23418 4059 23420
rect 4115 23418 4121 23420
rect 3875 23366 3877 23418
rect 4057 23366 4059 23418
rect 3813 23364 3819 23366
rect 3875 23364 3899 23366
rect 3955 23364 3979 23366
rect 4035 23364 4059 23366
rect 4115 23364 4121 23366
rect 3813 23355 4121 23364
rect 6104 23118 6132 24550
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6368 22976 6420 22982
rect 6368 22918 6420 22924
rect 4473 22876 4781 22885
rect 4473 22874 4479 22876
rect 4535 22874 4559 22876
rect 4615 22874 4639 22876
rect 4695 22874 4719 22876
rect 4775 22874 4781 22876
rect 4535 22822 4537 22874
rect 4717 22822 4719 22874
rect 4473 22820 4479 22822
rect 4535 22820 4559 22822
rect 4615 22820 4639 22822
rect 4695 22820 4719 22822
rect 4775 22820 4781 22822
rect 4473 22811 4781 22820
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 3813 22332 4121 22341
rect 3813 22330 3819 22332
rect 3875 22330 3899 22332
rect 3955 22330 3979 22332
rect 4035 22330 4059 22332
rect 4115 22330 4121 22332
rect 3875 22278 3877 22330
rect 4057 22278 4059 22330
rect 3813 22276 3819 22278
rect 3875 22276 3899 22278
rect 3955 22276 3979 22278
rect 4035 22276 4059 22278
rect 4115 22276 4121 22278
rect 3813 22267 4121 22276
rect 4473 21788 4781 21797
rect 4473 21786 4479 21788
rect 4535 21786 4559 21788
rect 4615 21786 4639 21788
rect 4695 21786 4719 21788
rect 4775 21786 4781 21788
rect 4535 21734 4537 21786
rect 4717 21734 4719 21786
rect 4473 21732 4479 21734
rect 4535 21732 4559 21734
rect 4615 21732 4639 21734
rect 4695 21732 4719 21734
rect 4775 21732 4781 21734
rect 4473 21723 4781 21732
rect 848 21548 900 21554
rect 848 21490 900 21496
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 860 21321 888 21490
rect 4344 21344 4396 21350
rect 846 21312 902 21321
rect 4344 21286 4396 21292
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 846 21247 902 21256
rect 3813 21244 4121 21253
rect 3813 21242 3819 21244
rect 3875 21242 3899 21244
rect 3955 21242 3979 21244
rect 4035 21242 4059 21244
rect 4115 21242 4121 21244
rect 3875 21190 3877 21242
rect 4057 21190 4059 21242
rect 3813 21188 3819 21190
rect 3875 21188 3899 21190
rect 3955 21188 3979 21190
rect 4035 21188 4059 21190
rect 4115 21188 4121 21190
rect 3813 21179 4121 21188
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20505 1440 20878
rect 3700 20800 3752 20806
rect 3700 20742 3752 20748
rect 1398 20496 1454 20505
rect 3712 20466 3740 20742
rect 1398 20431 1454 20440
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 846 19952 902 19961
rect 846 19887 902 19896
rect 860 19854 888 19887
rect 3436 19854 3464 20198
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3712 19310 3740 20402
rect 4356 20398 4384 21286
rect 4448 21010 4476 21286
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4540 20874 4568 21490
rect 5552 21486 5580 22510
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5920 21010 5948 22170
rect 6380 22030 6408 22918
rect 6748 22642 6776 24550
rect 7392 24206 7420 24550
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7392 23798 7420 24142
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8404 23866 8432 24006
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6472 21962 6500 22374
rect 6840 22234 6868 23122
rect 8312 22574 8340 23598
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6644 21956 6696 21962
rect 6644 21898 6696 21904
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 6012 20942 6040 21354
rect 6104 21010 6132 21422
rect 6472 21418 6500 21898
rect 6656 21486 6684 21898
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6460 21412 6512 21418
rect 6460 21354 6512 21360
rect 6840 21010 6868 21830
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 4528 20868 4580 20874
rect 4528 20810 4580 20816
rect 4473 20700 4781 20709
rect 4473 20698 4479 20700
rect 4535 20698 4559 20700
rect 4615 20698 4639 20700
rect 4695 20698 4719 20700
rect 4775 20698 4781 20700
rect 4535 20646 4537 20698
rect 4717 20646 4719 20698
rect 4473 20644 4479 20646
rect 4535 20644 4559 20646
rect 4615 20644 4639 20646
rect 4695 20644 4719 20646
rect 4775 20644 4781 20646
rect 4473 20635 4781 20644
rect 6380 20466 6408 20946
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 3813 20156 4121 20165
rect 3813 20154 3819 20156
rect 3875 20154 3899 20156
rect 3955 20154 3979 20156
rect 4035 20154 4059 20156
rect 4115 20154 4121 20156
rect 3875 20102 3877 20154
rect 4057 20102 4059 20154
rect 3813 20100 3819 20102
rect 3875 20100 3899 20102
rect 3955 20100 3979 20102
rect 4035 20100 4059 20102
rect 4115 20100 4121 20102
rect 3813 20091 4121 20100
rect 4264 19922 4292 20198
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 1400 19168 1452 19174
rect 1398 19136 1400 19145
rect 4160 19168 4212 19174
rect 1452 19136 1454 19145
rect 4160 19110 4212 19116
rect 1398 19071 1454 19080
rect 3813 19068 4121 19077
rect 3813 19066 3819 19068
rect 3875 19066 3899 19068
rect 3955 19066 3979 19068
rect 4035 19066 4059 19068
rect 4115 19066 4121 19068
rect 3875 19014 3877 19066
rect 4057 19014 4059 19066
rect 3813 19012 3819 19014
rect 3875 19012 3899 19014
rect 3955 19012 3979 19014
rect 4035 19012 4059 19014
rect 4115 19012 4121 19014
rect 3813 19003 4121 19012
rect 3976 18760 4028 18766
rect 4172 18748 4200 19110
rect 4264 18986 4292 19722
rect 4356 19378 4384 20334
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4448 19854 4476 20198
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4473 19612 4781 19621
rect 4473 19610 4479 19612
rect 4535 19610 4559 19612
rect 4615 19610 4639 19612
rect 4695 19610 4719 19612
rect 4775 19610 4781 19612
rect 4535 19558 4537 19610
rect 4717 19558 4719 19610
rect 4473 19556 4479 19558
rect 4535 19556 4559 19558
rect 4615 19556 4639 19558
rect 4695 19556 4719 19558
rect 4775 19556 4781 19558
rect 4473 19547 4781 19556
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4264 18958 4476 18986
rect 4448 18834 4476 18958
rect 4252 18828 4304 18834
rect 4436 18828 4488 18834
rect 4304 18788 4384 18816
rect 4252 18770 4304 18776
rect 4028 18720 4200 18748
rect 3976 18702 4028 18708
rect 848 18624 900 18630
rect 846 18592 848 18601
rect 900 18592 902 18601
rect 846 18527 902 18536
rect 3988 18222 4016 18702
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4264 18426 4292 18566
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4356 18358 4384 18788
rect 4436 18770 4488 18776
rect 4816 18766 4844 19654
rect 5092 18970 5120 19722
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4473 18524 4781 18533
rect 4473 18522 4479 18524
rect 4535 18522 4559 18524
rect 4615 18522 4639 18524
rect 4695 18522 4719 18524
rect 4775 18522 4781 18524
rect 4535 18470 4537 18522
rect 4717 18470 4719 18522
rect 4473 18468 4479 18470
rect 4535 18468 4559 18470
rect 4615 18468 4639 18470
rect 4695 18468 4719 18470
rect 4775 18468 4781 18470
rect 4473 18459 4781 18468
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 17785 1440 18022
rect 3813 17980 4121 17989
rect 3813 17978 3819 17980
rect 3875 17978 3899 17980
rect 3955 17978 3979 17980
rect 4035 17978 4059 17980
rect 4115 17978 4121 17980
rect 3875 17926 3877 17978
rect 4057 17926 4059 17978
rect 3813 17924 3819 17926
rect 3875 17924 3899 17926
rect 3955 17924 3979 17926
rect 4035 17924 4059 17926
rect 4115 17924 4121 17926
rect 3813 17915 4121 17924
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 846 17232 902 17241
rect 846 17167 848 17176
rect 900 17167 902 17176
rect 848 17138 900 17144
rect 3813 16892 4121 16901
rect 3813 16890 3819 16892
rect 3875 16890 3899 16892
rect 3955 16890 3979 16892
rect 4035 16890 4059 16892
rect 4115 16890 4121 16892
rect 3875 16838 3877 16890
rect 4057 16838 4059 16890
rect 3813 16836 3819 16838
rect 3875 16836 3899 16838
rect 3955 16836 3979 16838
rect 4035 16836 4059 16838
rect 4115 16836 4121 16838
rect 3813 16827 4121 16836
rect 848 16584 900 16590
rect 846 16552 848 16561
rect 900 16552 902 16561
rect 846 16487 902 16496
rect 4356 16250 4384 18294
rect 4908 17898 4936 18770
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18290 5028 18566
rect 5092 18426 5120 18702
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 5368 18222 5396 19926
rect 6380 19922 6408 20402
rect 6552 20324 6604 20330
rect 6552 20266 6604 20272
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6564 19854 6592 20266
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6656 18834 6684 19110
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6748 18766 6776 20742
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6932 19514 6960 19858
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7024 19310 7052 20946
rect 7300 20942 7328 21286
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7392 20874 7420 21286
rect 7380 20868 7432 20874
rect 7380 20810 7432 20816
rect 7472 20868 7524 20874
rect 7472 20810 7524 20816
rect 7484 20602 7512 20810
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7116 19514 7144 19790
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7208 18970 7236 19382
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 6736 18760 6788 18766
rect 6736 18702 6788 18708
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 4816 17870 4936 17898
rect 4816 17610 4844 17870
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4473 17436 4781 17445
rect 4473 17434 4479 17436
rect 4535 17434 4559 17436
rect 4615 17434 4639 17436
rect 4695 17434 4719 17436
rect 4775 17434 4781 17436
rect 4535 17382 4537 17434
rect 4717 17382 4719 17434
rect 4473 17380 4479 17382
rect 4535 17380 4559 17382
rect 4615 17380 4639 17382
rect 4695 17380 4719 17382
rect 4775 17380 4781 17382
rect 4473 17371 4781 17380
rect 4816 17134 4844 17546
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4908 16794 4936 17070
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4473 16348 4781 16357
rect 4473 16346 4479 16348
rect 4535 16346 4559 16348
rect 4615 16346 4639 16348
rect 4695 16346 4719 16348
rect 4775 16346 4781 16348
rect 4535 16294 4537 16346
rect 4717 16294 4719 16346
rect 4473 16292 4479 16294
rect 4535 16292 4559 16294
rect 4615 16292 4639 16294
rect 4695 16292 4719 16294
rect 4775 16292 4781 16294
rect 4473 16283 4781 16292
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 860 15881 888 16050
rect 846 15872 902 15881
rect 846 15807 902 15816
rect 3252 15706 3280 16050
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 3813 15804 4121 15813
rect 3813 15802 3819 15804
rect 3875 15802 3899 15804
rect 3955 15802 3979 15804
rect 4035 15802 4059 15804
rect 4115 15802 4121 15804
rect 3875 15750 3877 15802
rect 4057 15750 4059 15802
rect 3813 15748 3819 15750
rect 3875 15748 3899 15750
rect 3955 15748 3979 15750
rect 4035 15748 4059 15750
rect 4115 15748 4121 15750
rect 3813 15739 4121 15748
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 4264 15502 4292 15982
rect 5000 15706 5028 17138
rect 5368 16658 5396 18158
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6104 17882 6132 18090
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6288 17338 6316 17614
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6656 17270 6684 17478
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6840 17202 6868 17750
rect 7024 17338 7052 18634
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 17882 7144 18566
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 8220 17746 8248 19246
rect 8680 18426 8708 24754
rect 9048 24682 9076 26516
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9036 24676 9088 24682
rect 9036 24618 9088 24624
rect 8760 23656 8812 23662
rect 8760 23598 8812 23604
rect 8772 22234 8800 23598
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 8864 23118 8892 23462
rect 9048 23118 9076 23462
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 8864 22642 8892 23054
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 8864 22506 8892 22578
rect 9048 22574 9076 23054
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 8852 22500 8904 22506
rect 8852 22442 8904 22448
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8864 22166 8892 22442
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 8956 21554 8984 22374
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8944 21412 8996 21418
rect 8944 21354 8996 21360
rect 8956 20942 8984 21354
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 8772 19310 8800 19858
rect 8956 19514 8984 20198
rect 9048 19514 9076 22374
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8772 17814 8800 19246
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8956 18766 8984 19110
rect 9140 18970 9168 24754
rect 9692 24682 9720 26516
rect 10336 26466 10364 26516
rect 10428 26466 10456 26574
rect 10336 26438 10456 26466
rect 10200 25052 10508 25061
rect 10200 25050 10206 25052
rect 10262 25050 10286 25052
rect 10342 25050 10366 25052
rect 10422 25050 10446 25052
rect 10502 25050 10508 25052
rect 10262 24998 10264 25050
rect 10444 24998 10446 25050
rect 10200 24996 10206 24998
rect 10262 24996 10286 24998
rect 10342 24996 10366 24998
rect 10422 24996 10446 24998
rect 10502 24996 10508 24998
rect 10200 24987 10508 24996
rect 9864 24812 9916 24818
rect 9864 24754 9916 24760
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9324 23866 9352 24550
rect 9540 24508 9848 24517
rect 9540 24506 9546 24508
rect 9602 24506 9626 24508
rect 9682 24506 9706 24508
rect 9762 24506 9786 24508
rect 9842 24506 9848 24508
rect 9602 24454 9604 24506
rect 9784 24454 9786 24506
rect 9540 24452 9546 24454
rect 9602 24452 9626 24454
rect 9682 24452 9706 24454
rect 9762 24452 9786 24454
rect 9842 24452 9848 24454
rect 9540 24443 9848 24452
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9540 23420 9848 23429
rect 9540 23418 9546 23420
rect 9602 23418 9626 23420
rect 9682 23418 9706 23420
rect 9762 23418 9786 23420
rect 9842 23418 9848 23420
rect 9602 23366 9604 23418
rect 9784 23366 9786 23418
rect 9540 23364 9546 23366
rect 9602 23364 9626 23366
rect 9682 23364 9706 23366
rect 9762 23364 9786 23366
rect 9842 23364 9848 23366
rect 9540 23355 9848 23364
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9508 22778 9536 22918
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9220 22568 9272 22574
rect 9220 22510 9272 22516
rect 9232 22098 9260 22510
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9324 22114 9352 22374
rect 9416 22234 9444 22578
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9600 22438 9628 22510
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 9540 22332 9848 22341
rect 9540 22330 9546 22332
rect 9602 22330 9626 22332
rect 9682 22330 9706 22332
rect 9762 22330 9786 22332
rect 9842 22330 9848 22332
rect 9602 22278 9604 22330
rect 9784 22278 9786 22330
rect 9540 22276 9546 22278
rect 9602 22276 9626 22278
rect 9682 22276 9706 22278
rect 9762 22276 9786 22278
rect 9842 22276 9848 22278
rect 9540 22267 9848 22276
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9220 22092 9272 22098
rect 9324 22086 9444 22114
rect 9220 22034 9272 22040
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9232 21010 9260 21490
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 9416 20398 9444 22086
rect 9540 21244 9848 21253
rect 9540 21242 9546 21244
rect 9602 21242 9626 21244
rect 9682 21242 9706 21244
rect 9762 21242 9786 21244
rect 9842 21242 9848 21244
rect 9602 21190 9604 21242
rect 9784 21190 9786 21242
rect 9540 21188 9546 21190
rect 9602 21188 9626 21190
rect 9682 21188 9706 21190
rect 9762 21188 9786 21190
rect 9842 21188 9848 21190
rect 9540 21179 9848 21188
rect 9496 21004 9548 21010
rect 9496 20946 9548 20952
rect 9508 20602 9536 20946
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9416 19990 9444 20334
rect 9540 20156 9848 20165
rect 9540 20154 9546 20156
rect 9602 20154 9626 20156
rect 9682 20154 9706 20156
rect 9762 20154 9786 20156
rect 9842 20154 9848 20156
rect 9602 20102 9604 20154
rect 9784 20102 9786 20154
rect 9540 20100 9546 20102
rect 9602 20100 9626 20102
rect 9682 20100 9706 20102
rect 9762 20100 9786 20102
rect 9842 20100 9848 20102
rect 9540 20091 9848 20100
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9416 18766 9444 19654
rect 9540 19068 9848 19077
rect 9540 19066 9546 19068
rect 9602 19066 9626 19068
rect 9682 19066 9706 19068
rect 9762 19066 9786 19068
rect 9842 19066 9848 19068
rect 9602 19014 9604 19066
rect 9784 19014 9786 19066
rect 9540 19012 9546 19014
rect 9602 19012 9626 19014
rect 9682 19012 9706 19014
rect 9762 19012 9786 19014
rect 9842 19012 9848 19014
rect 9540 19003 9848 19012
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 8956 18154 8984 18702
rect 9416 18358 9444 18702
rect 9404 18352 9456 18358
rect 9404 18294 9456 18300
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16726 5488 16934
rect 7208 16794 7236 17478
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 5092 15706 5120 16118
rect 5184 16046 5212 16390
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 5368 15570 5396 16594
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 5460 15638 5488 16050
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 1412 15065 1440 15438
rect 3436 15366 3464 15438
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 3436 14958 3464 15302
rect 3620 15026 3648 15370
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3620 14618 3648 14962
rect 4264 14958 4292 15438
rect 6472 15434 6500 15846
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 15450 6684 15506
rect 6840 15502 6868 16050
rect 6932 15706 6960 16390
rect 7576 16250 7604 16390
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 6828 15496 6880 15502
rect 6656 15444 6828 15450
rect 6656 15438 6880 15444
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6656 15422 6868 15438
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4473 15260 4781 15269
rect 4473 15258 4479 15260
rect 4535 15258 4559 15260
rect 4615 15258 4639 15260
rect 4695 15258 4719 15260
rect 4775 15258 4781 15260
rect 4535 15206 4537 15258
rect 4717 15206 4719 15258
rect 4473 15204 4479 15206
rect 4535 15204 4559 15206
rect 4615 15204 4639 15206
rect 4695 15204 4719 15206
rect 4775 15204 4781 15206
rect 4473 15195 4781 15204
rect 4816 15162 4844 15302
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 3712 14618 3740 14894
rect 3813 14716 4121 14725
rect 3813 14714 3819 14716
rect 3875 14714 3899 14716
rect 3955 14714 3979 14716
rect 4035 14714 4059 14716
rect 4115 14714 4121 14716
rect 3875 14662 3877 14714
rect 4057 14662 4059 14714
rect 3813 14660 3819 14662
rect 3875 14660 3899 14662
rect 3955 14660 3979 14662
rect 4035 14660 4059 14662
rect 4115 14660 4121 14662
rect 3813 14651 4121 14660
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 846 14512 902 14521
rect 846 14447 902 14456
rect 5080 14476 5132 14482
rect 860 14414 888 14447
rect 5276 14464 5304 14962
rect 6656 14618 6684 15422
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 5132 14436 5304 14464
rect 5080 14418 5132 14424
rect 848 14408 900 14414
rect 848 14350 900 14356
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4356 14074 4384 14214
rect 4473 14172 4781 14181
rect 4473 14170 4479 14172
rect 4535 14170 4559 14172
rect 4615 14170 4639 14172
rect 4695 14170 4719 14172
rect 4775 14170 4781 14172
rect 4535 14118 4537 14170
rect 4717 14118 4719 14170
rect 4473 14116 4479 14118
rect 4535 14116 4559 14118
rect 4615 14116 4639 14118
rect 4695 14116 4719 14118
rect 4775 14116 4781 14118
rect 4473 14107 4781 14116
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 3813 13628 4121 13637
rect 3813 13626 3819 13628
rect 3875 13626 3899 13628
rect 3955 13626 3979 13628
rect 4035 13626 4059 13628
rect 4115 13626 4121 13628
rect 3875 13574 3877 13626
rect 4057 13574 4059 13626
rect 3813 13572 3819 13574
rect 3875 13572 3899 13574
rect 3955 13572 3979 13574
rect 4035 13572 4059 13574
rect 4115 13572 4121 13574
rect 3813 13563 4121 13572
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 13161 888 13262
rect 1584 13184 1636 13190
rect 846 13152 902 13161
rect 1584 13126 1636 13132
rect 846 13087 902 13096
rect 1596 12918 1624 13126
rect 4473 13084 4781 13093
rect 4473 13082 4479 13084
rect 4535 13082 4559 13084
rect 4615 13082 4639 13084
rect 4695 13082 4719 13084
rect 4775 13082 4781 13084
rect 4535 13030 4537 13082
rect 4717 13030 4719 13082
rect 4473 13028 4479 13030
rect 4535 13028 4559 13030
rect 4615 13028 4639 13030
rect 4695 13028 4719 13030
rect 4775 13028 4781 13030
rect 4473 13019 4781 13028
rect 1584 12912 1636 12918
rect 1584 12854 1636 12860
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 1412 12345 1440 12786
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 3813 12540 4121 12549
rect 3813 12538 3819 12540
rect 3875 12538 3899 12540
rect 3955 12538 3979 12540
rect 4035 12538 4059 12540
rect 4115 12538 4121 12540
rect 3875 12486 3877 12538
rect 4057 12486 4059 12538
rect 3813 12484 3819 12486
rect 3875 12484 3899 12486
rect 3955 12484 3979 12486
rect 4035 12484 4059 12486
rect 4115 12484 4121 12486
rect 3813 12475 4121 12484
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 846 11792 902 11801
rect 4356 11778 4384 12582
rect 4724 12306 4752 12650
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4816 12102 4844 12786
rect 5000 12220 5028 12786
rect 5276 12782 5304 14436
rect 7024 14414 7052 15574
rect 7300 15570 7328 16050
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7300 15162 7328 15506
rect 7392 15162 7420 15914
rect 8036 15706 8064 17478
rect 8220 16726 8248 17682
rect 8208 16720 8260 16726
rect 8772 16674 8800 17750
rect 9416 17678 9444 18158
rect 9540 17980 9848 17989
rect 9540 17978 9546 17980
rect 9602 17978 9626 17980
rect 9682 17978 9706 17980
rect 9762 17978 9786 17980
rect 9842 17978 9848 17980
rect 9602 17926 9604 17978
rect 9784 17926 9786 17978
rect 9540 17924 9546 17926
rect 9602 17924 9626 17926
rect 9682 17924 9706 17926
rect 9762 17924 9786 17926
rect 9842 17924 9848 17926
rect 9540 17915 9848 17924
rect 9876 17882 9904 24754
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9968 21622 9996 22374
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 10060 18970 10088 24754
rect 10612 24682 10640 26574
rect 10966 26516 11022 27316
rect 11610 26516 11666 27316
rect 12254 26516 12310 27316
rect 12898 26516 12954 27316
rect 13542 26516 13598 27316
rect 14186 26516 14242 27316
rect 14830 26516 14886 27316
rect 15474 26516 15530 27316
rect 16118 26516 16174 27316
rect 16762 26516 16818 27316
rect 17406 26516 17462 27316
rect 18050 26516 18106 27316
rect 20626 26516 20682 27316
rect 10980 24682 11008 26516
rect 11624 24818 11652 26516
rect 12268 24818 12296 26516
rect 12912 24818 12940 26516
rect 13556 24818 13584 26516
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 10600 24676 10652 24682
rect 10600 24618 10652 24624
rect 10968 24676 11020 24682
rect 10968 24618 11020 24624
rect 10200 23964 10508 23973
rect 10200 23962 10206 23964
rect 10262 23962 10286 23964
rect 10342 23962 10366 23964
rect 10422 23962 10446 23964
rect 10502 23962 10508 23964
rect 10262 23910 10264 23962
rect 10444 23910 10446 23962
rect 10200 23908 10206 23910
rect 10262 23908 10286 23910
rect 10342 23908 10366 23910
rect 10422 23908 10446 23910
rect 10502 23908 10508 23910
rect 10200 23899 10508 23908
rect 10200 22876 10508 22885
rect 10200 22874 10206 22876
rect 10262 22874 10286 22876
rect 10342 22874 10366 22876
rect 10422 22874 10446 22876
rect 10502 22874 10508 22876
rect 10262 22822 10264 22874
rect 10444 22822 10446 22874
rect 10200 22820 10206 22822
rect 10262 22820 10286 22822
rect 10342 22820 10366 22822
rect 10422 22820 10446 22822
rect 10502 22820 10508 22822
rect 10200 22811 10508 22820
rect 10200 21788 10508 21797
rect 10200 21786 10206 21788
rect 10262 21786 10286 21788
rect 10342 21786 10366 21788
rect 10422 21786 10446 21788
rect 10502 21786 10508 21788
rect 10262 21734 10264 21786
rect 10444 21734 10446 21786
rect 10200 21732 10206 21734
rect 10262 21732 10286 21734
rect 10342 21732 10366 21734
rect 10422 21732 10446 21734
rect 10502 21732 10508 21734
rect 10200 21723 10508 21732
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10336 21146 10364 21286
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10336 20942 10364 21082
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10200 20700 10508 20709
rect 10200 20698 10206 20700
rect 10262 20698 10286 20700
rect 10342 20698 10366 20700
rect 10422 20698 10446 20700
rect 10502 20698 10508 20700
rect 10262 20646 10264 20698
rect 10444 20646 10446 20698
rect 10200 20644 10206 20646
rect 10262 20644 10286 20646
rect 10342 20644 10366 20646
rect 10422 20644 10446 20646
rect 10502 20644 10508 20646
rect 10200 20635 10508 20644
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10612 19922 10640 20198
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10704 19786 10732 20946
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10200 19612 10508 19621
rect 10200 19610 10206 19612
rect 10262 19610 10286 19612
rect 10342 19610 10366 19612
rect 10422 19610 10446 19612
rect 10502 19610 10508 19612
rect 10262 19558 10264 19610
rect 10444 19558 10446 19610
rect 10200 19556 10206 19558
rect 10262 19556 10286 19558
rect 10342 19556 10366 19558
rect 10422 19556 10446 19558
rect 10502 19556 10508 19558
rect 10200 19547 10508 19556
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10200 18524 10508 18533
rect 10200 18522 10206 18524
rect 10262 18522 10286 18524
rect 10342 18522 10366 18524
rect 10422 18522 10446 18524
rect 10502 18522 10508 18524
rect 10262 18470 10264 18522
rect 10444 18470 10446 18522
rect 10200 18468 10206 18470
rect 10262 18468 10286 18470
rect 10342 18468 10366 18470
rect 10422 18468 10446 18470
rect 10502 18468 10508 18470
rect 10200 18459 10508 18468
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 11072 17814 11100 24754
rect 14200 24682 14228 26516
rect 14844 24818 14872 26516
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14188 24676 14240 24682
rect 14188 24618 14240 24624
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 11900 22778 11928 24550
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12360 23594 12388 23666
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 12360 22574 12388 23530
rect 12348 22568 12400 22574
rect 12348 22510 12400 22516
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11992 22094 12020 22374
rect 11992 22066 12112 22094
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11992 21554 12020 21830
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11256 21010 11284 21422
rect 12084 21418 12112 22066
rect 12544 22030 12572 24550
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11256 20874 11284 20946
rect 11808 20942 11836 21286
rect 11900 21010 11928 21286
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 12084 20874 12112 21354
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11440 19854 11468 20742
rect 12176 19922 12204 20946
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12636 20534 12664 20742
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 12176 18834 12204 19858
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 11532 17678 11560 18566
rect 11992 18290 12020 18566
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 9416 16794 9444 17614
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10200 17436 10508 17445
rect 10200 17434 10206 17436
rect 10262 17434 10286 17436
rect 10342 17434 10366 17436
rect 10422 17434 10446 17436
rect 10502 17434 10508 17436
rect 10262 17382 10264 17434
rect 10444 17382 10446 17434
rect 10200 17380 10206 17382
rect 10262 17380 10286 17382
rect 10342 17380 10366 17382
rect 10422 17380 10446 17382
rect 10502 17380 10508 17382
rect 10200 17371 10508 17380
rect 10796 17338 10824 17478
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 12176 17134 12204 18770
rect 12636 17882 12664 18770
rect 12728 18766 12756 20198
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 9540 16892 9848 16901
rect 9540 16890 9546 16892
rect 9602 16890 9626 16892
rect 9682 16890 9706 16892
rect 9762 16890 9786 16892
rect 9842 16890 9848 16892
rect 9602 16838 9604 16890
rect 9784 16838 9786 16890
rect 9540 16836 9546 16838
rect 9602 16836 9626 16838
rect 9682 16836 9706 16838
rect 9762 16836 9786 16838
rect 9842 16836 9848 16838
rect 9540 16827 9848 16836
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 11072 16726 11100 16934
rect 11060 16720 11112 16726
rect 8208 16662 8260 16668
rect 8588 16658 8892 16674
rect 11060 16662 11112 16668
rect 8588 16652 8904 16658
rect 8588 16646 8852 16652
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 7208 13802 7236 14418
rect 7392 14414 7420 15098
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7484 14618 7512 14894
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6932 12986 6960 13126
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 7024 12850 7052 13262
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 5276 12434 5304 12718
rect 6932 12442 6960 12718
rect 4908 12192 5028 12220
rect 5184 12406 5304 12434
rect 5356 12436 5408 12442
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4473 11996 4781 12005
rect 4473 11994 4479 11996
rect 4535 11994 4559 11996
rect 4615 11994 4639 11996
rect 4695 11994 4719 11996
rect 4775 11994 4781 11996
rect 4535 11942 4537 11994
rect 4717 11942 4719 11994
rect 4473 11940 4479 11942
rect 4535 11940 4559 11942
rect 4615 11940 4639 11942
rect 4695 11940 4719 11942
rect 4775 11940 4781 11942
rect 4473 11931 4781 11940
rect 4816 11898 4844 12038
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4172 11762 4384 11778
rect 846 11727 848 11736
rect 900 11727 902 11736
rect 4160 11756 4396 11762
rect 848 11698 900 11704
rect 4212 11750 4344 11756
rect 4160 11698 4212 11704
rect 4344 11698 4396 11704
rect 3813 11452 4121 11461
rect 3813 11450 3819 11452
rect 3875 11450 3899 11452
rect 3955 11450 3979 11452
rect 4035 11450 4059 11452
rect 4115 11450 4121 11452
rect 3875 11398 3877 11450
rect 4057 11398 4059 11450
rect 3813 11396 3819 11398
rect 3875 11396 3899 11398
rect 3955 11396 3979 11398
rect 4035 11396 4059 11398
rect 4115 11396 4121 11398
rect 3813 11387 4121 11396
rect 4356 11218 4384 11698
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4632 11150 4660 11494
rect 4908 11354 4936 12192
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 4473 10908 4781 10917
rect 4473 10906 4479 10908
rect 4535 10906 4559 10908
rect 4615 10906 4639 10908
rect 4695 10906 4719 10908
rect 4775 10906 4781 10908
rect 4535 10854 4537 10906
rect 4717 10854 4719 10906
rect 4473 10852 4479 10854
rect 4535 10852 4559 10854
rect 4615 10852 4639 10854
rect 4695 10852 4719 10854
rect 4775 10852 4781 10854
rect 4473 10843 4781 10852
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 848 10464 900 10470
rect 846 10432 848 10441
rect 900 10432 902 10441
rect 846 10367 902 10376
rect 3813 10364 4121 10373
rect 3813 10362 3819 10364
rect 3875 10362 3899 10364
rect 3955 10362 3979 10364
rect 4035 10362 4059 10364
rect 4115 10362 4121 10364
rect 3875 10310 3877 10362
rect 4057 10310 4059 10362
rect 3813 10308 3819 10310
rect 3875 10308 3899 10310
rect 3955 10308 3979 10310
rect 4035 10308 4059 10310
rect 4115 10308 4121 10310
rect 3813 10299 4121 10308
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 9625 1440 9862
rect 4473 9820 4781 9829
rect 4473 9818 4479 9820
rect 4535 9818 4559 9820
rect 4615 9818 4639 9820
rect 4695 9818 4719 9820
rect 4775 9818 4781 9820
rect 4535 9766 4537 9818
rect 4717 9766 4719 9818
rect 4473 9764 4479 9766
rect 4535 9764 4559 9766
rect 4615 9764 4639 9766
rect 4695 9764 4719 9766
rect 4775 9764 4781 9766
rect 4473 9755 4781 9764
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 4816 9382 4844 10610
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4908 9722 4936 9862
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5000 9654 5028 11494
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5092 10606 5120 11154
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 3813 9276 4121 9285
rect 3813 9274 3819 9276
rect 3875 9274 3899 9276
rect 3955 9274 3979 9276
rect 4035 9274 4059 9276
rect 4115 9274 4121 9276
rect 3875 9222 3877 9274
rect 4057 9222 4059 9274
rect 3813 9220 3819 9222
rect 3875 9220 3899 9222
rect 3955 9220 3979 9222
rect 4035 9220 4059 9222
rect 4115 9220 4121 9222
rect 3813 9211 4121 9220
rect 848 9104 900 9110
rect 846 9072 848 9081
rect 900 9072 902 9081
rect 846 9007 902 9016
rect 4473 8732 4781 8741
rect 4473 8730 4479 8732
rect 4535 8730 4559 8732
rect 4615 8730 4639 8732
rect 4695 8730 4719 8732
rect 4775 8730 4781 8732
rect 4535 8678 4537 8730
rect 4717 8678 4719 8730
rect 4473 8676 4479 8678
rect 4535 8676 4559 8678
rect 4615 8676 4639 8678
rect 4695 8676 4719 8678
rect 4775 8676 4781 8678
rect 4473 8667 4781 8676
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 3813 8188 4121 8197
rect 3813 8186 3819 8188
rect 3875 8186 3899 8188
rect 3955 8186 3979 8188
rect 4035 8186 4059 8188
rect 4115 8186 4121 8188
rect 3875 8134 3877 8186
rect 4057 8134 4059 8186
rect 3813 8132 3819 8134
rect 3875 8132 3899 8134
rect 3955 8132 3979 8134
rect 4035 8132 4059 8134
rect 4115 8132 4121 8134
rect 3813 8123 4121 8132
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 2596 7744 2648 7750
rect 846 7712 902 7721
rect 2596 7686 2648 7692
rect 846 7647 902 7656
rect 2608 7478 2636 7686
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6905 1440 7346
rect 4264 7342 4292 8230
rect 4356 7886 4384 8298
rect 4540 7954 4568 8366
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7546 4384 7822
rect 4540 7732 4568 7890
rect 4540 7704 4844 7732
rect 4473 7644 4781 7653
rect 4473 7642 4479 7644
rect 4535 7642 4559 7644
rect 4615 7642 4639 7644
rect 4695 7642 4719 7644
rect 4775 7642 4781 7644
rect 4535 7590 4537 7642
rect 4717 7590 4719 7642
rect 4473 7588 4479 7590
rect 4535 7588 4559 7590
rect 4615 7588 4639 7590
rect 4695 7588 4719 7590
rect 4775 7588 4781 7590
rect 4473 7579 4781 7588
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 3813 7100 4121 7109
rect 3813 7098 3819 7100
rect 3875 7098 3899 7100
rect 3955 7098 3979 7100
rect 4035 7098 4059 7100
rect 4115 7098 4121 7100
rect 3875 7046 3877 7098
rect 4057 7046 4059 7098
rect 3813 7044 3819 7046
rect 3875 7044 3899 7046
rect 3955 7044 3979 7046
rect 4035 7044 4059 7046
rect 4115 7044 4121 7046
rect 3813 7035 4121 7044
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 3813 6012 4121 6021
rect 3813 6010 3819 6012
rect 3875 6010 3899 6012
rect 3955 6010 3979 6012
rect 4035 6010 4059 6012
rect 4115 6010 4121 6012
rect 3875 5958 3877 6010
rect 4057 5958 4059 6010
rect 3813 5956 3819 5958
rect 3875 5956 3899 5958
rect 3955 5956 3979 5958
rect 4035 5956 4059 5958
rect 4115 5956 4121 5958
rect 3813 5947 4121 5956
rect 3813 4924 4121 4933
rect 3813 4922 3819 4924
rect 3875 4922 3899 4924
rect 3955 4922 3979 4924
rect 4035 4922 4059 4924
rect 4115 4922 4121 4924
rect 3875 4870 3877 4922
rect 4057 4870 4059 4922
rect 3813 4868 3819 4870
rect 3875 4868 3899 4870
rect 3955 4868 3979 4870
rect 4035 4868 4059 4870
rect 4115 4868 4121 4870
rect 3813 4859 4121 4868
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 4172 4146 4200 4490
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3813 3836 4121 3845
rect 3813 3834 3819 3836
rect 3875 3834 3899 3836
rect 3955 3834 3979 3836
rect 4035 3834 4059 3836
rect 4115 3834 4121 3836
rect 3875 3782 3877 3834
rect 4057 3782 4059 3834
rect 3813 3780 3819 3782
rect 3875 3780 3899 3782
rect 3955 3780 3979 3782
rect 4035 3780 4059 3782
rect 4115 3780 4121 3782
rect 3813 3771 4121 3780
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 3813 2748 4121 2757
rect 3813 2746 3819 2748
rect 3875 2746 3899 2748
rect 3955 2746 3979 2748
rect 4035 2746 4059 2748
rect 4115 2746 4121 2748
rect 3875 2694 3877 2746
rect 4057 2694 4059 2746
rect 3813 2692 3819 2694
rect 3875 2692 3899 2694
rect 3955 2692 3979 2694
rect 4035 2692 4059 2694
rect 4115 2692 4121 2694
rect 3813 2683 4121 2692
rect 4172 2650 4200 3062
rect 4264 2990 4292 7278
rect 4356 6934 4384 7482
rect 4816 7274 4844 7704
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 4816 6866 4844 7210
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4473 6556 4781 6565
rect 4473 6554 4479 6556
rect 4535 6554 4559 6556
rect 4615 6554 4639 6556
rect 4695 6554 4719 6556
rect 4775 6554 4781 6556
rect 4535 6502 4537 6554
rect 4717 6502 4719 6554
rect 4473 6500 4479 6502
rect 4535 6500 4559 6502
rect 4615 6500 4639 6502
rect 4695 6500 4719 6502
rect 4775 6500 4781 6502
rect 4473 6491 4781 6500
rect 4473 5468 4781 5477
rect 4473 5466 4479 5468
rect 4535 5466 4559 5468
rect 4615 5466 4639 5468
rect 4695 5466 4719 5468
rect 4775 5466 4781 5468
rect 4535 5414 4537 5466
rect 4717 5414 4719 5466
rect 4473 5412 4479 5414
rect 4535 5412 4559 5414
rect 4615 5412 4639 5414
rect 4695 5412 4719 5414
rect 4775 5412 4781 5414
rect 4473 5403 4781 5412
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4356 4282 4384 5170
rect 4473 4380 4781 4389
rect 4473 4378 4479 4380
rect 4535 4378 4559 4380
rect 4615 4378 4639 4380
rect 4695 4378 4719 4380
rect 4775 4378 4781 4380
rect 4535 4326 4537 4378
rect 4717 4326 4719 4378
rect 4473 4324 4479 4326
rect 4535 4324 4559 4326
rect 4615 4324 4639 4326
rect 4695 4324 4719 4326
rect 4775 4324 4781 4326
rect 4473 4315 4781 4324
rect 4816 4282 4844 5170
rect 4908 5166 4936 7890
rect 5000 6866 5028 9454
rect 5092 7954 5120 10066
rect 5184 8294 5212 12406
rect 5356 12378 5408 12384
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 10062 5304 10406
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5368 8106 5396 12378
rect 7116 12238 7144 12718
rect 7208 12434 7236 13738
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 7288 12436 7340 12442
rect 7208 12406 7288 12434
rect 7288 12378 7340 12384
rect 7392 12374 7420 12650
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7380 12368 7432 12374
rect 7432 12316 7512 12322
rect 7380 12310 7512 12316
rect 7392 12294 7512 12310
rect 8220 12306 8248 12582
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5460 11694 5488 11766
rect 5552 11694 5580 12038
rect 7116 11694 7144 12174
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11150 5856 11494
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5644 10810 5672 11018
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 8634 5488 10474
rect 7392 10062 7420 12038
rect 7484 11762 7512 12294
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 11830 8248 12242
rect 8312 12238 8340 12650
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11898 8524 12106
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11218 7696 11494
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7760 11150 7788 11562
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7852 10062 7880 11154
rect 8220 10130 8248 11766
rect 8588 11082 8616 16646
rect 8852 16594 8904 16600
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9784 15994 9812 16458
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9876 16250 9904 16390
rect 10060 16250 10088 16526
rect 10200 16348 10508 16357
rect 10200 16346 10206 16348
rect 10262 16346 10286 16348
rect 10342 16346 10366 16348
rect 10422 16346 10446 16348
rect 10502 16346 10508 16348
rect 10262 16294 10264 16346
rect 10444 16294 10446 16346
rect 10200 16292 10206 16294
rect 10262 16292 10286 16294
rect 10342 16292 10366 16294
rect 10422 16292 10446 16294
rect 10502 16292 10508 16294
rect 10200 16283 10508 16292
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9784 15966 9904 15994
rect 9540 15804 9848 15813
rect 9540 15802 9546 15804
rect 9602 15802 9626 15804
rect 9682 15802 9706 15804
rect 9762 15802 9786 15804
rect 9842 15802 9848 15804
rect 9602 15750 9604 15802
rect 9784 15750 9786 15802
rect 9540 15748 9546 15750
rect 9602 15748 9626 15750
rect 9682 15748 9706 15750
rect 9762 15748 9786 15750
rect 9842 15748 9848 15750
rect 9540 15739 9848 15748
rect 9876 15706 9904 15966
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8772 15162 8800 15506
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8680 12782 8708 15030
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9416 14618 9444 14962
rect 9540 14716 9848 14725
rect 9540 14714 9546 14716
rect 9602 14714 9626 14716
rect 9682 14714 9706 14716
rect 9762 14714 9786 14716
rect 9842 14714 9848 14716
rect 9602 14662 9604 14714
rect 9784 14662 9786 14714
rect 9540 14660 9546 14662
rect 9602 14660 9626 14662
rect 9682 14660 9706 14662
rect 9762 14660 9786 14662
rect 9842 14660 9848 14662
rect 9540 14651 9848 14660
rect 10060 14618 10088 16050
rect 11072 16046 11100 16662
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11072 15570 11100 15982
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10200 15260 10508 15269
rect 10200 15258 10206 15260
rect 10262 15258 10286 15260
rect 10342 15258 10366 15260
rect 10422 15258 10446 15260
rect 10502 15258 10508 15260
rect 10262 15206 10264 15258
rect 10444 15206 10446 15258
rect 10200 15204 10206 15206
rect 10262 15204 10286 15206
rect 10342 15204 10366 15206
rect 10422 15204 10446 15206
rect 10502 15204 10508 15206
rect 10200 15195 10508 15204
rect 10612 15162 10640 15302
rect 10704 15162 10732 15370
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 14346 9996 14418
rect 10244 14414 10272 14826
rect 10888 14822 10916 14894
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14618 10916 14758
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10692 14476 10744 14482
rect 10888 14464 10916 14554
rect 11072 14550 11100 15506
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10744 14436 10916 14464
rect 10692 14418 10744 14424
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9540 13628 9848 13637
rect 9540 13626 9546 13628
rect 9602 13626 9626 13628
rect 9682 13626 9706 13628
rect 9762 13626 9786 13628
rect 9842 13626 9848 13628
rect 9602 13574 9604 13626
rect 9784 13574 9786 13626
rect 9540 13572 9546 13574
rect 9602 13572 9626 13574
rect 9682 13572 9706 13574
rect 9762 13572 9786 13574
rect 9842 13572 9848 13574
rect 9540 13563 9848 13572
rect 9968 12986 9996 14282
rect 10200 14172 10508 14181
rect 10200 14170 10206 14172
rect 10262 14170 10286 14172
rect 10342 14170 10366 14172
rect 10422 14170 10446 14172
rect 10502 14170 10508 14172
rect 10262 14118 10264 14170
rect 10444 14118 10446 14170
rect 10200 14116 10206 14118
rect 10262 14116 10286 14118
rect 10342 14116 10366 14118
rect 10422 14116 10446 14118
rect 10502 14116 10508 14118
rect 10200 14107 10508 14116
rect 10200 13084 10508 13093
rect 10200 13082 10206 13084
rect 10262 13082 10286 13084
rect 10342 13082 10366 13084
rect 10422 13082 10446 13084
rect 10502 13082 10508 13084
rect 10262 13030 10264 13082
rect 10444 13030 10446 13082
rect 10200 13028 10206 13030
rect 10262 13028 10286 13030
rect 10342 13028 10366 13030
rect 10422 13028 10446 13030
rect 10502 13028 10508 13030
rect 10200 13019 10508 13028
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 9540 12540 9848 12549
rect 9540 12538 9546 12540
rect 9602 12538 9626 12540
rect 9682 12538 9706 12540
rect 9762 12538 9786 12540
rect 9842 12538 9848 12540
rect 9602 12486 9604 12538
rect 9784 12486 9786 12538
rect 9540 12484 9546 12486
rect 9602 12484 9626 12486
rect 9682 12484 9706 12486
rect 9762 12484 9786 12486
rect 9842 12484 9848 12486
rect 9540 12475 9848 12484
rect 10428 12442 10456 12786
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 10060 11898 10088 12106
rect 10200 11996 10508 12005
rect 10200 11994 10206 11996
rect 10262 11994 10286 11996
rect 10342 11994 10366 11996
rect 10422 11994 10446 11996
rect 10502 11994 10508 11996
rect 10262 11942 10264 11994
rect 10444 11942 10446 11994
rect 10200 11940 10206 11942
rect 10262 11940 10286 11942
rect 10342 11940 10366 11942
rect 10422 11940 10446 11942
rect 10502 11940 10508 11942
rect 10200 11931 10508 11940
rect 10612 11898 10640 12174
rect 10888 11898 10916 12786
rect 11072 12646 11100 14486
rect 11808 14278 11836 17002
rect 12084 16794 12112 17070
rect 12360 17066 12388 17546
rect 12636 17202 12664 17614
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12360 16590 12388 17002
rect 12636 16794 12664 17138
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 15026 11928 16390
rect 12360 16250 12388 16526
rect 12728 16250 12756 17138
rect 12820 16590 12848 24550
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13096 20466 13124 20742
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13280 18358 13308 18566
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13096 17882 13124 18226
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12912 16250 12940 16934
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14414 11928 14962
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12360 14618 12388 14826
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12452 14482 12480 15030
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14482 12848 14758
rect 13004 14482 13032 15982
rect 13096 15094 13124 16594
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11808 13938 11836 14214
rect 11992 14074 12020 14214
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 13004 13802 13032 14418
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 13004 13394 13032 13738
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9540 11452 9848 11461
rect 9540 11450 9546 11452
rect 9602 11450 9626 11452
rect 9682 11450 9706 11452
rect 9762 11450 9786 11452
rect 9842 11450 9848 11452
rect 9602 11398 9604 11450
rect 9784 11398 9786 11450
rect 9540 11396 9546 11398
rect 9602 11396 9626 11398
rect 9682 11396 9706 11398
rect 9762 11396 9786 11398
rect 9842 11396 9848 11398
rect 9540 11387 9848 11396
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8588 10198 8616 11018
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7300 9722 7328 9862
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7392 9654 7420 9862
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5368 8078 5488 8106
rect 5644 8090 5672 8434
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5092 7834 5120 7890
rect 5092 7806 5304 7834
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5092 7546 5120 7686
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7002 5212 7686
rect 5276 7274 5304 7806
rect 5368 7410 5396 7890
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 5000 6254 5028 6802
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 5778 5028 6190
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5092 5370 5120 5510
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4908 4690 4936 5102
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 5184 4486 5212 5510
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4816 3466 4844 3946
rect 4908 3942 4936 4082
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3534 4936 3878
rect 5000 3738 5028 4422
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4473 3292 4781 3301
rect 4473 3290 4479 3292
rect 4535 3290 4559 3292
rect 4615 3290 4639 3292
rect 4695 3290 4719 3292
rect 4775 3290 4781 3292
rect 4535 3238 4537 3290
rect 4717 3238 4719 3290
rect 4473 3236 4479 3238
rect 4535 3236 4559 3238
rect 4615 3236 4639 3238
rect 4695 3236 4719 3238
rect 4775 3236 4781 3238
rect 4473 3227 4781 3236
rect 4816 3194 4844 3402
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4540 2650 4568 2994
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4540 2446 4568 2586
rect 4724 2514 4752 2790
rect 4908 2650 4936 3470
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5276 2514 5304 6938
rect 5368 5302 5396 7346
rect 5460 7206 5488 8078
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 5736 7342 5764 7822
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 5460 7002 5488 7142
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 7024 6798 7052 7142
rect 7116 6798 7144 7754
rect 7300 7546 7328 7822
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7392 6798 7420 9318
rect 8036 9178 8064 9454
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7484 7002 7512 7346
rect 8220 7342 8248 10066
rect 8588 9178 8616 10134
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8588 9042 8616 9114
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5370 5580 5646
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5460 4826 5488 5170
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5644 4078 5672 4558
rect 5828 4146 5856 4626
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 3194 6960 3470
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 2582 6868 2790
rect 6932 2650 6960 2994
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 7024 2446 7052 6598
rect 7392 5914 7420 6734
rect 7944 6118 7972 7278
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7300 4146 7328 4694
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7484 4282 7512 4490
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7300 3534 7328 4082
rect 7576 4078 7604 4490
rect 7668 4078 7696 5102
rect 7944 4162 7972 6054
rect 7852 4134 7972 4162
rect 7852 4078 7880 4134
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7576 3618 7604 4014
rect 7944 3738 7972 4014
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7576 3590 7696 3618
rect 7668 3534 7696 3590
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 3194 7696 3470
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7116 2650 7144 2926
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7208 2514 7236 2926
rect 7288 2576 7340 2582
rect 7392 2564 7420 3130
rect 7340 2536 7420 2564
rect 7288 2518 7340 2524
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 8036 2446 8064 7142
rect 8404 6798 8432 7142
rect 8588 6866 8616 8978
rect 9324 7410 9352 11222
rect 10060 11218 10088 11494
rect 10520 11354 10548 11630
rect 11072 11354 11100 12582
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11440 11218 11468 12038
rect 11624 11694 11652 12106
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11900 11626 11928 12106
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11532 11150 11560 11494
rect 11900 11354 11928 11562
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 10200 10908 10508 10917
rect 10200 10906 10206 10908
rect 10262 10906 10286 10908
rect 10342 10906 10366 10908
rect 10422 10906 10446 10908
rect 10502 10906 10508 10908
rect 10262 10854 10264 10906
rect 10444 10854 10446 10906
rect 10200 10852 10206 10854
rect 10262 10852 10286 10854
rect 10342 10852 10366 10854
rect 10422 10852 10446 10854
rect 10502 10852 10508 10854
rect 10200 10843 10508 10852
rect 9540 10364 9848 10373
rect 9540 10362 9546 10364
rect 9602 10362 9626 10364
rect 9682 10362 9706 10364
rect 9762 10362 9786 10364
rect 9842 10362 9848 10364
rect 9602 10310 9604 10362
rect 9784 10310 9786 10362
rect 9540 10308 9546 10310
rect 9602 10308 9626 10310
rect 9682 10308 9706 10310
rect 9762 10308 9786 10310
rect 9842 10308 9848 10310
rect 9540 10299 9848 10308
rect 10200 9820 10508 9829
rect 10200 9818 10206 9820
rect 10262 9818 10286 9820
rect 10342 9818 10366 9820
rect 10422 9818 10446 9820
rect 10502 9818 10508 9820
rect 10262 9766 10264 9818
rect 10444 9766 10446 9818
rect 10200 9764 10206 9766
rect 10262 9764 10286 9766
rect 10342 9764 10366 9766
rect 10422 9764 10446 9766
rect 10502 9764 10508 9766
rect 10200 9755 10508 9764
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9416 8974 9444 9318
rect 9540 9276 9848 9285
rect 9540 9274 9546 9276
rect 9602 9274 9626 9276
rect 9682 9274 9706 9276
rect 9762 9274 9786 9276
rect 9842 9274 9848 9276
rect 9602 9222 9604 9274
rect 9784 9222 9786 9274
rect 9540 9220 9546 9222
rect 9602 9220 9626 9222
rect 9682 9220 9706 9222
rect 9762 9220 9786 9222
rect 9842 9220 9848 9222
rect 9540 9211 9848 9220
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 10612 8906 10640 9522
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10200 8732 10508 8741
rect 10200 8730 10206 8732
rect 10262 8730 10286 8732
rect 10342 8730 10366 8732
rect 10422 8730 10446 8732
rect 10502 8730 10508 8732
rect 10262 8678 10264 8730
rect 10444 8678 10446 8730
rect 10200 8676 10206 8678
rect 10262 8676 10286 8678
rect 10342 8676 10366 8678
rect 10422 8676 10446 8678
rect 10502 8676 10508 8678
rect 10200 8667 10508 8676
rect 10612 8548 10640 8842
rect 10704 8838 10732 9454
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10520 8520 10640 8548
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 9540 8188 9848 8197
rect 9540 8186 9546 8188
rect 9602 8186 9626 8188
rect 9682 8186 9706 8188
rect 9762 8186 9786 8188
rect 9842 8186 9848 8188
rect 9602 8134 9604 8186
rect 9784 8134 9786 8186
rect 9540 8132 9546 8134
rect 9602 8132 9626 8134
rect 9682 8132 9706 8134
rect 9762 8132 9786 8134
rect 9842 8132 9848 8134
rect 9540 8123 9848 8132
rect 10060 8022 10088 8434
rect 10244 8090 10272 8434
rect 10520 8294 10548 8520
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10520 7954 10548 8230
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10200 7644 10508 7653
rect 10200 7642 10206 7644
rect 10262 7642 10286 7644
rect 10342 7642 10366 7644
rect 10422 7642 10446 7644
rect 10502 7642 10508 7644
rect 10262 7590 10264 7642
rect 10444 7590 10446 7642
rect 10200 7588 10206 7590
rect 10262 7588 10286 7590
rect 10342 7588 10366 7590
rect 10422 7588 10446 7590
rect 10502 7588 10508 7590
rect 10200 7579 10508 7588
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8588 6746 8616 6802
rect 8772 6798 8800 7278
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 8760 6792 8812 6798
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8312 5166 8340 6190
rect 8404 6186 8432 6734
rect 8588 6718 8708 6746
rect 8760 6734 8812 6740
rect 8576 6656 8628 6662
rect 8680 6644 8708 6718
rect 8680 6616 8800 6644
rect 8576 6598 8628 6604
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4282 8156 4422
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8496 4010 8524 6258
rect 8588 5114 8616 6598
rect 8772 6390 8800 6616
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8680 5914 8708 6190
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8588 5086 8708 5114
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4690 8616 4966
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8680 2446 8708 5086
rect 9324 2446 9352 7142
rect 9540 7100 9848 7109
rect 9540 7098 9546 7100
rect 9602 7098 9626 7100
rect 9682 7098 9706 7100
rect 9762 7098 9786 7100
rect 9842 7098 9848 7100
rect 9602 7046 9604 7098
rect 9784 7046 9786 7098
rect 9540 7044 9546 7046
rect 9602 7044 9626 7046
rect 9682 7044 9706 7046
rect 9762 7044 9786 7046
rect 9842 7044 9848 7046
rect 9540 7035 9848 7044
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9600 6458 9628 6734
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9540 6012 9848 6021
rect 9540 6010 9546 6012
rect 9602 6010 9626 6012
rect 9682 6010 9706 6012
rect 9762 6010 9786 6012
rect 9842 6010 9848 6012
rect 9602 5958 9604 6010
rect 9784 5958 9786 6010
rect 9540 5956 9546 5958
rect 9602 5956 9626 5958
rect 9682 5956 9706 5958
rect 9762 5956 9786 5958
rect 9842 5956 9848 5958
rect 9540 5947 9848 5956
rect 9540 4924 9848 4933
rect 9540 4922 9546 4924
rect 9602 4922 9626 4924
rect 9682 4922 9706 4924
rect 9762 4922 9786 4924
rect 9842 4922 9848 4924
rect 9602 4870 9604 4922
rect 9784 4870 9786 4922
rect 9540 4868 9546 4870
rect 9602 4868 9626 4870
rect 9682 4868 9706 4870
rect 9762 4868 9786 4870
rect 9842 4868 9848 4870
rect 9540 4859 9848 4868
rect 9540 3836 9848 3845
rect 9540 3834 9546 3836
rect 9602 3834 9626 3836
rect 9682 3834 9706 3836
rect 9762 3834 9786 3836
rect 9842 3834 9848 3836
rect 9602 3782 9604 3834
rect 9784 3782 9786 3834
rect 9540 3780 9546 3782
rect 9602 3780 9626 3782
rect 9682 3780 9706 3782
rect 9762 3780 9786 3782
rect 9842 3780 9848 3782
rect 9540 3771 9848 3780
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9876 3058 9904 3402
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9540 2748 9848 2757
rect 9540 2746 9546 2748
rect 9602 2746 9626 2748
rect 9682 2746 9706 2748
rect 9762 2746 9786 2748
rect 9842 2746 9848 2748
rect 9602 2694 9604 2746
rect 9784 2694 9786 2746
rect 9540 2692 9546 2694
rect 9602 2692 9626 2694
rect 9682 2692 9706 2694
rect 9762 2692 9786 2694
rect 9842 2692 9848 2694
rect 9540 2683 9848 2692
rect 9968 2446 9996 6598
rect 10200 6556 10508 6565
rect 10200 6554 10206 6556
rect 10262 6554 10286 6556
rect 10342 6554 10366 6556
rect 10422 6554 10446 6556
rect 10502 6554 10508 6556
rect 10262 6502 10264 6554
rect 10444 6502 10446 6554
rect 10200 6500 10206 6502
rect 10262 6500 10286 6502
rect 10342 6500 10366 6502
rect 10422 6500 10446 6502
rect 10502 6500 10508 6502
rect 10200 6491 10508 6500
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 4010 10088 6258
rect 10612 5710 10640 8298
rect 10704 7886 10732 8774
rect 10796 8498 10824 9522
rect 10876 9512 10928 9518
rect 10928 9460 11008 9466
rect 10876 9454 11008 9460
rect 10888 9438 11008 9454
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 8634 10916 9318
rect 10980 9178 11008 9438
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11152 8968 11204 8974
rect 10980 8916 11152 8922
rect 10980 8910 11204 8916
rect 10980 8906 11192 8910
rect 10968 8900 11192 8906
rect 11020 8894 11192 8900
rect 10968 8842 11020 8848
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10200 5468 10508 5477
rect 10200 5466 10206 5468
rect 10262 5466 10286 5468
rect 10342 5466 10366 5468
rect 10422 5466 10446 5468
rect 10502 5466 10508 5468
rect 10262 5414 10264 5466
rect 10444 5414 10446 5466
rect 10200 5412 10206 5414
rect 10262 5412 10286 5414
rect 10342 5412 10366 5414
rect 10422 5412 10446 5414
rect 10502 5412 10508 5414
rect 10200 5403 10508 5412
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 10200 4380 10508 4389
rect 10200 4378 10206 4380
rect 10262 4378 10286 4380
rect 10342 4378 10366 4380
rect 10422 4378 10446 4380
rect 10502 4378 10508 4380
rect 10262 4326 10264 4378
rect 10444 4326 10446 4378
rect 10200 4324 10206 4326
rect 10262 4324 10286 4326
rect 10342 4324 10366 4326
rect 10422 4324 10446 4326
rect 10502 4324 10508 4326
rect 10200 4315 10508 4324
rect 10612 4214 10640 4490
rect 10704 4298 10732 6394
rect 10796 4570 10824 8434
rect 10980 6914 11008 8842
rect 11256 8650 11284 9386
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11164 8622 11284 8650
rect 11164 8430 11192 8622
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11164 7954 11192 8366
rect 11256 7954 11284 8434
rect 11992 8430 12020 8774
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12360 8362 12388 11222
rect 12452 11218 12480 12038
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12636 11082 12664 12174
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 11694 12848 11834
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 10888 6886 11008 6914
rect 10888 6458 10916 6886
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10980 6458 11008 6734
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10888 5914 10916 6258
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10888 4826 10916 5714
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11152 4616 11204 4622
rect 10796 4542 11100 4570
rect 11152 4558 11204 4564
rect 10704 4270 10824 4298
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10612 3738 10640 4150
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10704 3738 10732 4082
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10060 3194 10088 3334
rect 10200 3292 10508 3301
rect 10200 3290 10206 3292
rect 10262 3290 10286 3292
rect 10342 3290 10366 3292
rect 10422 3290 10446 3292
rect 10502 3290 10508 3292
rect 10262 3238 10264 3290
rect 10444 3238 10446 3290
rect 10200 3236 10206 3238
rect 10262 3236 10286 3238
rect 10342 3236 10366 3238
rect 10422 3236 10446 3238
rect 10502 3236 10508 3238
rect 10200 3227 10508 3236
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 3252 800 3280 2382
rect 3896 800 3924 2382
rect 4356 1306 4384 2382
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 4473 2204 4781 2213
rect 4473 2202 4479 2204
rect 4535 2202 4559 2204
rect 4615 2202 4639 2204
rect 4695 2202 4719 2204
rect 4775 2202 4781 2204
rect 4535 2150 4537 2202
rect 4717 2150 4719 2202
rect 4473 2148 4479 2150
rect 4535 2148 4559 2150
rect 4615 2148 4639 2150
rect 4695 2148 4719 2150
rect 4775 2148 4781 2150
rect 4473 2139 4781 2148
rect 4356 1278 4568 1306
rect 4540 800 4568 1278
rect 5184 800 5212 2314
rect 5828 800 5856 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 800 6500 2246
rect 7116 800 7144 2382
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 9048 800 9076 2246
rect 9692 800 9720 2246
rect 10200 2204 10508 2213
rect 10200 2202 10206 2204
rect 10262 2202 10286 2204
rect 10342 2202 10366 2204
rect 10422 2202 10446 2204
rect 10502 2202 10508 2204
rect 10262 2150 10264 2202
rect 10444 2150 10446 2202
rect 10200 2148 10206 2150
rect 10262 2148 10286 2150
rect 10342 2148 10366 2150
rect 10422 2148 10446 2150
rect 10502 2148 10508 2150
rect 10200 2139 10508 2148
rect 10336 870 10456 898
rect 10336 800 10364 870
rect 18 0 74 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10428 762 10456 870
rect 10612 762 10640 2382
rect 10796 2378 10824 4270
rect 11072 3924 11100 4542
rect 11164 4282 11192 4558
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 10980 3896 11100 3924
rect 10980 2650 11008 3896
rect 11164 3602 11192 4218
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11256 2650 11284 7890
rect 12360 6914 12388 8298
rect 12360 6886 12572 6914
rect 12544 6254 12572 6886
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 5302 11560 5510
rect 11520 5296 11572 5302
rect 11520 5238 11572 5244
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11348 4826 11376 5170
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 12544 3670 12572 6190
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11900 2650 11928 3334
rect 12084 3126 12112 3538
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12636 2650 12664 11018
rect 12820 9110 12848 11630
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12728 5914 12756 6190
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 13096 2774 13124 11562
rect 13188 10674 13216 18022
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13280 11218 13308 13330
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13556 10742 13584 17206
rect 13648 17202 13676 24550
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14292 22574 14320 23462
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 20602 14228 21830
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14108 19854 14136 20198
rect 14476 20058 14504 24754
rect 15488 24682 15516 26516
rect 16132 25650 16160 26516
rect 16132 25622 16344 25650
rect 15927 25052 16235 25061
rect 15927 25050 15933 25052
rect 15989 25050 16013 25052
rect 16069 25050 16093 25052
rect 16149 25050 16173 25052
rect 16229 25050 16235 25052
rect 15989 24998 15991 25050
rect 16171 24998 16173 25050
rect 15927 24996 15933 24998
rect 15989 24996 16013 24998
rect 16069 24996 16093 24998
rect 16149 24996 16173 24998
rect 16229 24996 16235 24998
rect 15927 24987 16235 24996
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15476 24676 15528 24682
rect 15476 24618 15528 24624
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14936 23866 14964 24550
rect 15267 24508 15575 24517
rect 15267 24506 15273 24508
rect 15329 24506 15353 24508
rect 15409 24506 15433 24508
rect 15489 24506 15513 24508
rect 15569 24506 15575 24508
rect 15329 24454 15331 24506
rect 15511 24454 15513 24506
rect 15267 24452 15273 24454
rect 15329 24452 15353 24454
rect 15409 24452 15433 24454
rect 15489 24452 15513 24454
rect 15569 24452 15575 24454
rect 15267 24443 15575 24452
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15580 23866 15608 24006
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14752 23322 14780 23598
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14936 23118 14964 23802
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 14924 23112 14976 23118
rect 14924 23054 14976 23060
rect 15028 22710 15056 23462
rect 15267 23420 15575 23429
rect 15267 23418 15273 23420
rect 15329 23418 15353 23420
rect 15409 23418 15433 23420
rect 15489 23418 15513 23420
rect 15569 23418 15575 23420
rect 15329 23366 15331 23418
rect 15511 23366 15513 23418
rect 15267 23364 15273 23366
rect 15329 23364 15353 23366
rect 15409 23364 15433 23366
rect 15489 23364 15513 23366
rect 15569 23364 15575 23366
rect 15267 23355 15575 23364
rect 15672 23186 15700 23598
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14660 22030 14688 22374
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14752 21894 14780 22374
rect 14936 22030 14964 22510
rect 15028 22216 15056 22646
rect 15267 22332 15575 22341
rect 15267 22330 15273 22332
rect 15329 22330 15353 22332
rect 15409 22330 15433 22332
rect 15489 22330 15513 22332
rect 15569 22330 15575 22332
rect 15329 22278 15331 22330
rect 15511 22278 15513 22330
rect 15267 22276 15273 22278
rect 15329 22276 15353 22278
rect 15409 22276 15433 22278
rect 15489 22276 15513 22278
rect 15569 22276 15575 22278
rect 15267 22267 15575 22276
rect 15672 22234 15700 23122
rect 15660 22228 15712 22234
rect 15028 22188 15148 22216
rect 15120 22098 15148 22188
rect 15660 22170 15712 22176
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14936 21418 14964 21966
rect 14924 21412 14976 21418
rect 14924 21354 14976 21360
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14660 19922 14688 20878
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 14752 19854 14780 20946
rect 15028 20942 15056 22034
rect 15120 21622 15148 22034
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15120 21146 15148 21422
rect 15267 21244 15575 21253
rect 15267 21242 15273 21244
rect 15329 21242 15353 21244
rect 15409 21242 15433 21244
rect 15489 21242 15513 21244
rect 15569 21242 15575 21244
rect 15329 21190 15331 21242
rect 15511 21190 15513 21242
rect 15267 21188 15273 21190
rect 15329 21188 15353 21190
rect 15409 21188 15433 21190
rect 15489 21188 15513 21190
rect 15569 21188 15575 21190
rect 15267 21179 15575 21188
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14108 18902 14136 19790
rect 14752 18902 14780 19790
rect 14844 19378 14872 20402
rect 14936 20058 14964 20402
rect 15267 20156 15575 20165
rect 15267 20154 15273 20156
rect 15329 20154 15353 20156
rect 15409 20154 15433 20156
rect 15489 20154 15513 20156
rect 15569 20154 15575 20156
rect 15329 20102 15331 20154
rect 15511 20102 15513 20154
rect 15267 20100 15273 20102
rect 15329 20100 15353 20102
rect 15409 20100 15433 20102
rect 15489 20100 15513 20102
rect 15569 20100 15575 20102
rect 15267 20091 15575 20100
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13740 16046 13768 17070
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13832 13870 13860 14350
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13530 13860 13806
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 11898 13860 12718
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13740 10810 13860 10826
rect 13728 10804 13860 10810
rect 13780 10798 13860 10804
rect 13728 10746 13780 10752
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13188 6798 13216 7754
rect 13280 7546 13308 10610
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13556 10266 13584 10542
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13740 9654 13768 10610
rect 13832 9654 13860 10798
rect 14016 10674 14044 18566
rect 14108 16114 14136 18634
rect 14568 18426 14596 18634
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14752 17882 14780 18158
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14108 15706 14136 16050
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14844 15570 14872 19314
rect 15267 19068 15575 19077
rect 15267 19066 15273 19068
rect 15329 19066 15353 19068
rect 15409 19066 15433 19068
rect 15489 19066 15513 19068
rect 15569 19066 15575 19068
rect 15329 19014 15331 19066
rect 15511 19014 15513 19066
rect 15267 19012 15273 19014
rect 15329 19012 15353 19014
rect 15409 19012 15433 19014
rect 15489 19012 15513 19014
rect 15569 19012 15575 19014
rect 15267 19003 15575 19012
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15304 18426 15332 18634
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 15267 17980 15575 17989
rect 15267 17978 15273 17980
rect 15329 17978 15353 17980
rect 15409 17978 15433 17980
rect 15489 17978 15513 17980
rect 15569 17978 15575 17980
rect 15329 17926 15331 17978
rect 15511 17926 15513 17978
rect 15267 17924 15273 17926
rect 15329 17924 15353 17926
rect 15409 17924 15433 17926
rect 15489 17924 15513 17926
rect 15569 17924 15575 17926
rect 15267 17915 15575 17924
rect 15672 17746 15700 18090
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 17338 15240 17614
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15267 16892 15575 16901
rect 15267 16890 15273 16892
rect 15329 16890 15353 16892
rect 15409 16890 15433 16892
rect 15489 16890 15513 16892
rect 15569 16890 15575 16892
rect 15329 16838 15331 16890
rect 15511 16838 15513 16890
rect 15267 16836 15273 16838
rect 15329 16836 15353 16838
rect 15409 16836 15433 16838
rect 15489 16836 15513 16838
rect 15569 16836 15575 16838
rect 15267 16827 15575 16836
rect 15764 16250 15792 24754
rect 16316 24682 16344 25622
rect 16776 24818 16804 26516
rect 17420 24818 17448 26516
rect 18064 24818 18092 26516
rect 20640 24818 20668 26516
rect 21654 25052 21962 25061
rect 21654 25050 21660 25052
rect 21716 25050 21740 25052
rect 21796 25050 21820 25052
rect 21876 25050 21900 25052
rect 21956 25050 21962 25052
rect 21716 24998 21718 25050
rect 21898 24998 21900 25050
rect 21654 24996 21660 24998
rect 21716 24996 21740 24998
rect 21796 24996 21820 24998
rect 21876 24996 21900 24998
rect 21956 24996 21962 24998
rect 21654 24987 21962 24996
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 23664 24812 23716 24818
rect 23664 24754 23716 24760
rect 16304 24676 16356 24682
rect 16304 24618 16356 24624
rect 15927 23964 16235 23973
rect 15927 23962 15933 23964
rect 15989 23962 16013 23964
rect 16069 23962 16093 23964
rect 16149 23962 16173 23964
rect 16229 23962 16235 23964
rect 15989 23910 15991 23962
rect 16171 23910 16173 23962
rect 15927 23908 15933 23910
rect 15989 23908 16013 23910
rect 16069 23908 16093 23910
rect 16149 23908 16173 23910
rect 16229 23908 16235 23910
rect 15927 23899 16235 23908
rect 15927 22876 16235 22885
rect 15927 22874 15933 22876
rect 15989 22874 16013 22876
rect 16069 22874 16093 22876
rect 16149 22874 16173 22876
rect 16229 22874 16235 22876
rect 15989 22822 15991 22874
rect 16171 22822 16173 22874
rect 15927 22820 15933 22822
rect 15989 22820 16013 22822
rect 16069 22820 16093 22822
rect 16149 22820 16173 22822
rect 16229 22820 16235 22822
rect 15927 22811 16235 22820
rect 15927 21788 16235 21797
rect 15927 21786 15933 21788
rect 15989 21786 16013 21788
rect 16069 21786 16093 21788
rect 16149 21786 16173 21788
rect 16229 21786 16235 21788
rect 15989 21734 15991 21786
rect 16171 21734 16173 21786
rect 15927 21732 15933 21734
rect 15989 21732 16013 21734
rect 16069 21732 16093 21734
rect 16149 21732 16173 21734
rect 16229 21732 16235 21734
rect 15927 21723 16235 21732
rect 15927 20700 16235 20709
rect 15927 20698 15933 20700
rect 15989 20698 16013 20700
rect 16069 20698 16093 20700
rect 16149 20698 16173 20700
rect 16229 20698 16235 20700
rect 15989 20646 15991 20698
rect 16171 20646 16173 20698
rect 15927 20644 15933 20646
rect 15989 20644 16013 20646
rect 16069 20644 16093 20646
rect 16149 20644 16173 20646
rect 16229 20644 16235 20646
rect 15927 20635 16235 20644
rect 16408 20058 16436 24754
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 16868 24206 16896 24550
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16868 23798 16896 24142
rect 17604 23866 17632 24550
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 16856 23792 16908 23798
rect 16856 23734 16908 23740
rect 18340 23730 18368 24550
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17052 22574 17080 23462
rect 18064 23118 18092 23462
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18340 23050 18368 23666
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 18328 23044 18380 23050
rect 18328 22986 18380 22992
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17420 22642 17448 22918
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 17040 22568 17092 22574
rect 17040 22510 17092 22516
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 16580 22160 16632 22166
rect 16580 22102 16632 22108
rect 16592 22030 16620 22102
rect 16684 22098 16712 22442
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16776 21962 16804 22510
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 17236 22030 17264 22374
rect 17420 22234 17448 22578
rect 20640 22574 20668 23598
rect 20916 22778 20944 24550
rect 20994 24508 21302 24517
rect 20994 24506 21000 24508
rect 21056 24506 21080 24508
rect 21136 24506 21160 24508
rect 21216 24506 21240 24508
rect 21296 24506 21302 24508
rect 21056 24454 21058 24506
rect 21238 24454 21240 24506
rect 20994 24452 21000 24454
rect 21056 24452 21080 24454
rect 21136 24452 21160 24454
rect 21216 24452 21240 24454
rect 21296 24452 21302 24454
rect 20994 24443 21302 24452
rect 21654 23964 21962 23973
rect 21654 23962 21660 23964
rect 21716 23962 21740 23964
rect 21796 23962 21820 23964
rect 21876 23962 21900 23964
rect 21956 23962 21962 23964
rect 21716 23910 21718 23962
rect 21898 23910 21900 23962
rect 21654 23908 21660 23910
rect 21716 23908 21740 23910
rect 21796 23908 21820 23910
rect 21876 23908 21900 23910
rect 21956 23908 21962 23910
rect 21654 23899 21962 23908
rect 20994 23420 21302 23429
rect 20994 23418 21000 23420
rect 21056 23418 21080 23420
rect 21136 23418 21160 23420
rect 21216 23418 21240 23420
rect 21296 23418 21302 23420
rect 21056 23366 21058 23418
rect 21238 23366 21240 23418
rect 20994 23364 21000 23366
rect 21056 23364 21080 23366
rect 21136 23364 21160 23366
rect 21216 23364 21240 23366
rect 21296 23364 21302 23366
rect 20994 23355 21302 23364
rect 22756 23186 22784 24686
rect 23676 24585 23704 24754
rect 23662 24576 23718 24585
rect 23662 24511 23718 24520
rect 23020 24268 23072 24274
rect 23020 24210 23072 24216
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 21654 22876 21962 22885
rect 21654 22874 21660 22876
rect 21716 22874 21740 22876
rect 21796 22874 21820 22876
rect 21876 22874 21900 22876
rect 21956 22874 21962 22876
rect 21716 22822 21718 22874
rect 21898 22822 21900 22874
rect 21654 22820 21660 22822
rect 21716 22820 21740 22822
rect 21796 22820 21820 22822
rect 21876 22820 21900 22822
rect 21956 22820 21962 22822
rect 21654 22811 21962 22820
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 17500 22500 17552 22506
rect 17500 22442 17552 22448
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16684 19854 16712 21830
rect 16776 21486 16804 21898
rect 17420 21554 17448 22170
rect 17512 22098 17540 22442
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 17592 22092 17644 22098
rect 17592 22034 17644 22040
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16960 20942 16988 21286
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 17328 20602 17356 20946
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 17512 20398 17540 22034
rect 17604 21010 17632 22034
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 17788 21486 17816 21966
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 18064 21146 18092 21490
rect 20916 21486 20944 22374
rect 20994 22332 21302 22341
rect 20994 22330 21000 22332
rect 21056 22330 21080 22332
rect 21136 22330 21160 22332
rect 21216 22330 21240 22332
rect 21296 22330 21302 22332
rect 21056 22278 21058 22330
rect 21238 22278 21240 22330
rect 20994 22276 21000 22278
rect 21056 22276 21080 22278
rect 21136 22276 21160 22278
rect 21216 22276 21240 22278
rect 21296 22276 21302 22278
rect 20994 22267 21302 22276
rect 21654 21788 21962 21797
rect 21654 21786 21660 21788
rect 21716 21786 21740 21788
rect 21796 21786 21820 21788
rect 21876 21786 21900 21788
rect 21956 21786 21962 21788
rect 21716 21734 21718 21786
rect 21898 21734 21900 21786
rect 21654 21732 21660 21734
rect 21716 21732 21740 21734
rect 21796 21732 21820 21734
rect 21876 21732 21900 21734
rect 21956 21732 21962 21734
rect 21654 21723 21962 21732
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 18144 21072 18196 21078
rect 18144 21014 18196 21020
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17868 20392 17920 20398
rect 18156 20346 18184 21014
rect 19812 20942 19840 21286
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19444 20602 19472 20742
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19536 20534 19564 20742
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19904 20398 19932 21422
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20548 20534 20576 21286
rect 20732 20942 20760 21422
rect 20812 21412 20864 21418
rect 20812 21354 20864 21360
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 20602 20760 20742
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 20824 20466 20852 21354
rect 20916 21078 20944 21422
rect 20994 21244 21302 21253
rect 20994 21242 21000 21244
rect 21056 21242 21080 21244
rect 21136 21242 21160 21244
rect 21216 21242 21240 21244
rect 21296 21242 21302 21244
rect 21056 21190 21058 21242
rect 21238 21190 21240 21242
rect 20994 21188 21000 21190
rect 21056 21188 21080 21190
rect 21136 21188 21160 21190
rect 21216 21188 21240 21190
rect 21296 21188 21302 21190
rect 20994 21179 21302 21188
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 20916 20534 20944 21014
rect 22756 21010 22784 23122
rect 23032 22574 23060 24210
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23676 23905 23704 24142
rect 23662 23896 23718 23905
rect 23662 23831 23718 23840
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23400 23225 23428 23666
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 23386 23216 23442 23225
rect 23386 23151 23442 23160
rect 23664 22636 23716 22642
rect 23664 22578 23716 22584
rect 23020 22568 23072 22574
rect 23676 22545 23704 22578
rect 23020 22510 23072 22516
rect 23662 22536 23718 22545
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21284 20806 21312 20878
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 21284 20466 21312 20742
rect 21654 20700 21962 20709
rect 21654 20698 21660 20700
rect 21716 20698 21740 20700
rect 21796 20698 21820 20700
rect 21876 20698 21900 20700
rect 21956 20698 21962 20700
rect 21716 20646 21718 20698
rect 21898 20646 21900 20698
rect 21654 20644 21660 20646
rect 21716 20644 21740 20646
rect 21796 20644 21820 20646
rect 21876 20644 21900 20646
rect 21956 20644 21962 20646
rect 21654 20635 21962 20644
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 17920 20340 18184 20346
rect 17868 20334 18184 20340
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 17880 20318 18184 20334
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 19922 16804 20198
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 15856 19718 15884 19790
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15856 18970 15884 19654
rect 15927 19612 16235 19621
rect 15927 19610 15933 19612
rect 15989 19610 16013 19612
rect 16069 19610 16093 19612
rect 16149 19610 16173 19612
rect 16229 19610 16235 19612
rect 15989 19558 15991 19610
rect 16171 19558 16173 19610
rect 15927 19556 15933 19558
rect 15989 19556 16013 19558
rect 16069 19556 16093 19558
rect 16149 19556 16173 19558
rect 16229 19556 16235 19558
rect 15927 19547 16235 19556
rect 16960 19378 16988 19858
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15927 18524 16235 18533
rect 15927 18522 15933 18524
rect 15989 18522 16013 18524
rect 16069 18522 16093 18524
rect 16149 18522 16173 18524
rect 16229 18522 16235 18524
rect 15989 18470 15991 18522
rect 16171 18470 16173 18522
rect 15927 18468 15933 18470
rect 15989 18468 16013 18470
rect 16069 18468 16093 18470
rect 16149 18468 16173 18470
rect 16229 18468 16235 18470
rect 15927 18459 16235 18468
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15856 18086 15884 18226
rect 16960 18222 16988 19314
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 18064 18426 18092 18702
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 15856 17678 15884 18022
rect 16592 17746 16620 18022
rect 17328 17882 17356 18226
rect 18156 18222 18184 20318
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18800 19514 18828 19790
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18984 19378 19012 20198
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 17880 17678 17908 18022
rect 18156 17814 18184 18158
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 15856 16794 15884 17614
rect 15927 17436 16235 17445
rect 15927 17434 15933 17436
rect 15989 17434 16013 17436
rect 16069 17434 16093 17436
rect 16149 17434 16173 17436
rect 16229 17434 16235 17436
rect 15989 17382 15991 17434
rect 16171 17382 16173 17434
rect 15927 17380 15933 17382
rect 15989 17380 16013 17382
rect 16069 17380 16093 17382
rect 16149 17380 16173 17382
rect 16229 17380 16235 17382
rect 15927 17371 16235 17380
rect 17880 17270 17908 17614
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15948 16658 15976 16934
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 16132 16590 16160 17002
rect 16224 16726 16252 17070
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 15927 16348 16235 16357
rect 15927 16346 15933 16348
rect 15989 16346 16013 16348
rect 16069 16346 16093 16348
rect 16149 16346 16173 16348
rect 16229 16346 16235 16348
rect 15989 16294 15991 16346
rect 16171 16294 16173 16346
rect 15927 16292 15933 16294
rect 15989 16292 16013 16294
rect 16069 16292 16093 16294
rect 16149 16292 16173 16294
rect 16229 16292 16235 16294
rect 15927 16283 16235 16292
rect 17972 16250 18000 16390
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 15267 15804 15575 15813
rect 15267 15802 15273 15804
rect 15329 15802 15353 15804
rect 15409 15802 15433 15804
rect 15489 15802 15513 15804
rect 15569 15802 15575 15804
rect 15329 15750 15331 15802
rect 15511 15750 15513 15802
rect 15267 15748 15273 15750
rect 15329 15748 15353 15750
rect 15409 15748 15433 15750
rect 15489 15748 15513 15750
rect 15569 15748 15575 15750
rect 15267 15739 15575 15748
rect 17972 15586 18000 15982
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 17880 15558 18000 15586
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14476 14618 14504 15302
rect 15212 14770 15240 15302
rect 15672 15026 15700 15506
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 15927 15260 16235 15269
rect 15927 15258 15933 15260
rect 15989 15258 16013 15260
rect 16069 15258 16093 15260
rect 16149 15258 16173 15260
rect 16229 15258 16235 15260
rect 15989 15206 15991 15258
rect 16171 15206 16173 15258
rect 15927 15204 15933 15206
rect 15989 15204 16013 15206
rect 16069 15204 16093 15206
rect 16149 15204 16173 15206
rect 16229 15204 16235 15206
rect 15927 15195 16235 15204
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15120 14742 15240 14770
rect 15120 14618 15148 14742
rect 15267 14716 15575 14725
rect 15267 14714 15273 14716
rect 15329 14714 15353 14716
rect 15409 14714 15433 14716
rect 15489 14714 15513 14716
rect 15569 14714 15575 14716
rect 15329 14662 15331 14714
rect 15511 14662 15513 14714
rect 15267 14660 15273 14662
rect 15329 14660 15353 14662
rect 15409 14660 15433 14662
rect 15489 14660 15513 14662
rect 15569 14660 15575 14662
rect 15267 14651 15575 14660
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15672 14550 15700 14962
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 14108 13870 14136 14282
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14476 14074 14504 14214
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 15580 13938 15608 14418
rect 17144 14414 17172 15302
rect 17880 15026 17908 15558
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 15094 18000 15438
rect 18064 15162 18092 16390
rect 18156 16046 18184 17750
rect 18248 17202 18276 19314
rect 19812 18834 19840 20334
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19260 18222 19288 18702
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19536 18426 19564 18566
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19812 18154 19840 18770
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19996 18426 20024 18702
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20916 18290 20944 20198
rect 20994 20156 21302 20165
rect 20994 20154 21000 20156
rect 21056 20154 21080 20156
rect 21136 20154 21160 20156
rect 21216 20154 21240 20156
rect 21296 20154 21302 20156
rect 21056 20102 21058 20154
rect 21238 20102 21240 20154
rect 20994 20100 21000 20102
rect 21056 20100 21080 20102
rect 21136 20100 21160 20102
rect 21216 20100 21240 20102
rect 21296 20100 21302 20102
rect 20994 20091 21302 20100
rect 21654 19612 21962 19621
rect 21654 19610 21660 19612
rect 21716 19610 21740 19612
rect 21796 19610 21820 19612
rect 21876 19610 21900 19612
rect 21956 19610 21962 19612
rect 21716 19558 21718 19610
rect 21898 19558 21900 19610
rect 21654 19556 21660 19558
rect 21716 19556 21740 19558
rect 21796 19556 21820 19558
rect 21876 19556 21900 19558
rect 21956 19556 21962 19558
rect 21654 19547 21962 19556
rect 20994 19068 21302 19077
rect 20994 19066 21000 19068
rect 21056 19066 21080 19068
rect 21136 19066 21160 19068
rect 21216 19066 21240 19068
rect 21296 19066 21302 19068
rect 21056 19014 21058 19066
rect 21238 19014 21240 19066
rect 20994 19012 21000 19014
rect 21056 19012 21080 19014
rect 21136 19012 21160 19014
rect 21216 19012 21240 19014
rect 21296 19012 21302 19014
rect 20994 19003 21302 19012
rect 22100 18692 22152 18698
rect 22100 18634 22152 18640
rect 21654 18524 21962 18533
rect 21654 18522 21660 18524
rect 21716 18522 21740 18524
rect 21796 18522 21820 18524
rect 21876 18522 21900 18524
rect 21956 18522 21962 18524
rect 21716 18470 21718 18522
rect 21898 18470 21900 18522
rect 21654 18468 21660 18470
rect 21716 18468 21740 18470
rect 21796 18468 21820 18470
rect 21876 18468 21900 18470
rect 21956 18468 21962 18470
rect 21654 18459 21962 18468
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17328 14414 17356 14758
rect 17604 14414 17632 14826
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15672 13870 15700 14350
rect 15927 14172 16235 14181
rect 15927 14170 15933 14172
rect 15989 14170 16013 14172
rect 16069 14170 16093 14172
rect 16149 14170 16173 14172
rect 16229 14170 16235 14172
rect 15989 14118 15991 14170
rect 16171 14118 16173 14170
rect 15927 14116 15933 14118
rect 15989 14116 16013 14118
rect 16069 14116 16093 14118
rect 16149 14116 16173 14118
rect 16229 14116 16235 14118
rect 15927 14107 16235 14116
rect 17604 14074 17632 14350
rect 17880 14278 17908 14826
rect 17972 14618 18000 15030
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17880 13938 17908 14214
rect 18064 14074 18092 14962
rect 18248 14770 18276 16934
rect 18340 16794 18368 17138
rect 19536 16794 19564 17138
rect 18328 16788 18380 16794
rect 19524 16788 19576 16794
rect 18380 16748 18460 16776
rect 18328 16730 18380 16736
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18156 14742 18276 14770
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 14108 13394 14136 13806
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 15267 13628 15575 13637
rect 15267 13626 15273 13628
rect 15329 13626 15353 13628
rect 15409 13626 15433 13628
rect 15489 13626 15513 13628
rect 15569 13626 15575 13628
rect 15329 13574 15331 13626
rect 15511 13574 15513 13626
rect 15267 13572 15273 13574
rect 15329 13572 15353 13574
rect 15409 13572 15433 13574
rect 15489 13572 15513 13574
rect 15569 13572 15575 13574
rect 15267 13563 15575 13572
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14108 12986 14136 13330
rect 15764 13326 15792 13670
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14292 10198 14320 10406
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13372 9178 13400 9454
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13280 6254 13308 6802
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13280 5778 13308 6190
rect 13372 6118 13400 8774
rect 13464 8634 13492 9522
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 9042 13952 9318
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13740 8430 13768 8910
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13648 8090 13676 8366
rect 13924 8090 13952 8434
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14660 7954 14688 9046
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 13556 6934 13584 7890
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14476 7410 14504 7754
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7546 14596 7686
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13464 5710 13492 6598
rect 13556 6458 13584 6870
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13832 5574 13860 6258
rect 14292 5846 14320 6326
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13740 2922 13768 3606
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13096 2746 13400 2774
rect 13372 2650 13400 2746
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13832 2446 13860 5510
rect 14292 2650 14320 5782
rect 14384 5778 14412 6190
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14384 5370 14412 5714
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14568 4826 14596 5170
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14660 3058 14688 7890
rect 14936 5370 14964 12786
rect 15267 12540 15575 12549
rect 15267 12538 15273 12540
rect 15329 12538 15353 12540
rect 15409 12538 15433 12540
rect 15489 12538 15513 12540
rect 15569 12538 15575 12540
rect 15329 12486 15331 12538
rect 15511 12486 15513 12538
rect 15267 12484 15273 12486
rect 15329 12484 15353 12486
rect 15409 12484 15433 12486
rect 15489 12484 15513 12486
rect 15569 12484 15575 12486
rect 15267 12475 15575 12484
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15580 11762 15608 12242
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11762 15792 12174
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15580 11642 15608 11698
rect 15580 11614 15700 11642
rect 15267 11452 15575 11461
rect 15267 11450 15273 11452
rect 15329 11450 15353 11452
rect 15409 11450 15433 11452
rect 15489 11450 15513 11452
rect 15569 11450 15575 11452
rect 15329 11398 15331 11450
rect 15511 11398 15513 11450
rect 15267 11396 15273 11398
rect 15329 11396 15353 11398
rect 15409 11396 15433 11398
rect 15489 11396 15513 11398
rect 15569 11396 15575 11398
rect 15267 11387 15575 11396
rect 15672 11354 15700 11614
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15304 10742 15332 11290
rect 15764 10742 15792 11698
rect 15856 11642 15884 13126
rect 15927 13084 16235 13093
rect 15927 13082 15933 13084
rect 15989 13082 16013 13084
rect 16069 13082 16093 13084
rect 16149 13082 16173 13084
rect 16229 13082 16235 13084
rect 15989 13030 15991 13082
rect 16171 13030 16173 13082
rect 15927 13028 15933 13030
rect 15989 13028 16013 13030
rect 16069 13028 16093 13030
rect 16149 13028 16173 13030
rect 16229 13028 16235 13030
rect 15927 13019 16235 13028
rect 17052 12714 17080 13670
rect 17144 13530 17172 13806
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17236 13326 17264 13738
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 15927 11996 16235 12005
rect 15927 11994 15933 11996
rect 15989 11994 16013 11996
rect 16069 11994 16093 11996
rect 16149 11994 16173 11996
rect 16229 11994 16235 11996
rect 15989 11942 15991 11994
rect 16171 11942 16173 11994
rect 15927 11940 15933 11942
rect 15989 11940 16013 11942
rect 16069 11940 16093 11942
rect 16149 11940 16173 11942
rect 16229 11940 16235 11942
rect 15927 11931 16235 11940
rect 15856 11626 16068 11642
rect 15856 11620 16080 11626
rect 15856 11614 16028 11620
rect 15856 11150 15884 11614
rect 16028 11562 16080 11568
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 15948 11218 15976 11494
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15927 10908 16235 10917
rect 15927 10906 15933 10908
rect 15989 10906 16013 10908
rect 16069 10906 16093 10908
rect 16149 10906 16173 10908
rect 16229 10906 16235 10908
rect 15989 10854 15991 10906
rect 16171 10854 16173 10906
rect 15927 10852 15933 10854
rect 15989 10852 16013 10854
rect 16069 10852 16093 10854
rect 16149 10852 16173 10854
rect 16229 10852 16235 10854
rect 15927 10843 16235 10852
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15267 10364 15575 10373
rect 15267 10362 15273 10364
rect 15329 10362 15353 10364
rect 15409 10362 15433 10364
rect 15489 10362 15513 10364
rect 15569 10362 15575 10364
rect 15329 10310 15331 10362
rect 15511 10310 15513 10362
rect 15267 10308 15273 10310
rect 15329 10308 15353 10310
rect 15409 10308 15433 10310
rect 15489 10308 15513 10310
rect 15569 10308 15575 10310
rect 15267 10299 15575 10308
rect 15856 10130 15884 10406
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15948 10010 15976 10474
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16132 10062 16160 10406
rect 15856 9982 15976 10010
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9722 15424 9862
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15267 9276 15575 9285
rect 15267 9274 15273 9276
rect 15329 9274 15353 9276
rect 15409 9274 15433 9276
rect 15489 9274 15513 9276
rect 15569 9274 15575 9276
rect 15329 9222 15331 9274
rect 15511 9222 15513 9274
rect 15267 9220 15273 9222
rect 15329 9220 15353 9222
rect 15409 9220 15433 9222
rect 15489 9220 15513 9222
rect 15569 9220 15575 9222
rect 15267 9211 15575 9220
rect 15672 8498 15700 9318
rect 15764 9178 15792 9454
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15267 8188 15575 8197
rect 15267 8186 15273 8188
rect 15329 8186 15353 8188
rect 15409 8186 15433 8188
rect 15489 8186 15513 8188
rect 15569 8186 15575 8188
rect 15329 8134 15331 8186
rect 15511 8134 15513 8186
rect 15267 8132 15273 8134
rect 15329 8132 15353 8134
rect 15409 8132 15433 8134
rect 15489 8132 15513 8134
rect 15569 8132 15575 8134
rect 15267 8123 15575 8132
rect 15672 8022 15700 8434
rect 15856 8090 15884 9982
rect 15927 9820 16235 9829
rect 15927 9818 15933 9820
rect 15989 9818 16013 9820
rect 16069 9818 16093 9820
rect 16149 9818 16173 9820
rect 16229 9818 16235 9820
rect 15989 9766 15991 9818
rect 16171 9766 16173 9818
rect 15927 9764 15933 9766
rect 15989 9764 16013 9766
rect 16069 9764 16093 9766
rect 16149 9764 16173 9766
rect 16229 9764 16235 9766
rect 15927 9755 16235 9764
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 9042 16252 9318
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16316 8906 16344 11154
rect 16408 11150 16436 11494
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16500 11082 16528 12242
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17052 11830 17080 12174
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17144 11898 17172 12038
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9042 16436 10066
rect 17696 10062 17724 10950
rect 18156 10266 18184 14742
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18248 11150 18276 12582
rect 18340 11218 18368 16594
rect 18432 16590 18460 16748
rect 19524 16730 19576 16736
rect 19812 16658 19840 18090
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 20994 17980 21302 17989
rect 20994 17978 21000 17980
rect 21056 17978 21080 17980
rect 21136 17978 21160 17980
rect 21216 17978 21240 17980
rect 21296 17978 21302 17980
rect 21056 17926 21058 17978
rect 21238 17926 21240 17978
rect 20994 17924 21000 17926
rect 21056 17924 21080 17926
rect 21136 17924 21160 17926
rect 21216 17924 21240 17926
rect 21296 17924 21302 17926
rect 20994 17915 21302 17924
rect 21376 17678 21404 18022
rect 22112 17882 22140 18634
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21654 17436 21962 17445
rect 21654 17434 21660 17436
rect 21716 17434 21740 17436
rect 21796 17434 21820 17436
rect 21876 17434 21900 17436
rect 21956 17434 21962 17436
rect 21716 17382 21718 17434
rect 21898 17382 21900 17434
rect 21654 17380 21660 17382
rect 21716 17380 21740 17382
rect 21796 17380 21820 17382
rect 21876 17380 21900 17382
rect 21956 17380 21962 17382
rect 21654 17371 21962 17380
rect 20994 16892 21302 16901
rect 20994 16890 21000 16892
rect 21056 16890 21080 16892
rect 21136 16890 21160 16892
rect 21216 16890 21240 16892
rect 21296 16890 21302 16892
rect 21056 16838 21058 16890
rect 21238 16838 21240 16890
rect 20994 16836 21000 16838
rect 21056 16836 21080 16838
rect 21136 16836 21160 16838
rect 21216 16836 21240 16838
rect 21296 16836 21302 16838
rect 20994 16827 21302 16836
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 20720 16584 20772 16590
rect 22020 16561 22048 16662
rect 20720 16526 20772 16532
rect 22006 16552 22062 16561
rect 18800 16250 18828 16526
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 14958 18552 16050
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18892 15026 18920 15506
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18432 14618 18460 14894
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 19076 12782 19104 15982
rect 19904 15706 19932 16390
rect 19996 16250 20024 16390
rect 20732 16250 20760 16526
rect 22006 16487 22062 16496
rect 21654 16348 21962 16357
rect 21654 16346 21660 16348
rect 21716 16346 21740 16348
rect 21796 16346 21820 16348
rect 21876 16346 21900 16348
rect 21956 16346 21962 16348
rect 21716 16294 21718 16346
rect 21898 16294 21900 16346
rect 21654 16292 21660 16294
rect 21716 16292 21740 16294
rect 21796 16292 21820 16294
rect 21876 16292 21900 16294
rect 21956 16292 21962 16294
rect 21654 16283 21962 16292
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 22204 16114 22232 17750
rect 22296 17678 22324 18090
rect 22388 17882 22416 18566
rect 22572 18290 22600 18566
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22572 17814 22600 18226
rect 22756 18222 22784 20946
rect 23032 18834 23060 22510
rect 23662 22471 23718 22480
rect 23112 22432 23164 22438
rect 23112 22374 23164 22380
rect 23124 20942 23152 22374
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23572 21888 23624 21894
rect 23676 21865 23704 21966
rect 23572 21830 23624 21836
rect 23662 21856 23718 21865
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23400 20505 23428 20878
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23386 20496 23442 20505
rect 23386 20431 23442 20440
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23216 18970 23244 19314
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 22560 17808 22612 17814
rect 22560 17750 22612 17756
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 20994 15804 21302 15813
rect 20994 15802 21000 15804
rect 21056 15802 21080 15804
rect 21136 15802 21160 15804
rect 21216 15802 21240 15804
rect 21296 15802 21302 15804
rect 21056 15750 21058 15802
rect 21238 15750 21240 15802
rect 20994 15748 21000 15750
rect 21056 15748 21080 15750
rect 21136 15748 21160 15750
rect 21216 15748 21240 15750
rect 21296 15748 21302 15750
rect 20994 15739 21302 15748
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 21560 15570 21588 15982
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 22020 15502 22048 15982
rect 22204 15638 22232 16050
rect 22192 15632 22244 15638
rect 22192 15574 22244 15580
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21376 15162 21404 15302
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 20994 14716 21302 14725
rect 20994 14714 21000 14716
rect 21056 14714 21080 14716
rect 21136 14714 21160 14716
rect 21216 14714 21240 14716
rect 21296 14714 21302 14716
rect 21056 14662 21058 14714
rect 21238 14662 21240 14714
rect 20994 14660 21000 14662
rect 21056 14660 21080 14662
rect 21136 14660 21160 14662
rect 21216 14660 21240 14662
rect 21296 14660 21302 14662
rect 20994 14651 21302 14660
rect 21468 14618 21496 15302
rect 21560 15094 21588 15302
rect 21654 15260 21962 15269
rect 21654 15258 21660 15260
rect 21716 15258 21740 15260
rect 21796 15258 21820 15260
rect 21876 15258 21900 15260
rect 21956 15258 21962 15260
rect 21716 15206 21718 15258
rect 21898 15206 21900 15258
rect 21654 15204 21660 15206
rect 21716 15204 21740 15206
rect 21796 15204 21820 15206
rect 21876 15204 21900 15206
rect 21956 15204 21962 15206
rect 21654 15195 21962 15204
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21652 14618 21680 14962
rect 22020 14958 22048 15438
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 22112 14414 22140 14894
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14550 22324 14758
rect 22284 14544 22336 14550
rect 22284 14486 22336 14492
rect 23124 14482 23152 18158
rect 23216 16574 23244 18770
rect 23308 18465 23336 19314
rect 23400 19145 23428 19450
rect 23386 19136 23442 19145
rect 23386 19071 23442 19080
rect 23492 18766 23520 20742
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23294 18456 23350 18465
rect 23294 18391 23350 18400
rect 23584 18290 23612 21830
rect 23662 21791 23718 21800
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 21185 23704 21286
rect 23662 21176 23718 21185
rect 23662 21111 23718 21120
rect 23662 19816 23718 19825
rect 23662 19751 23718 19760
rect 23676 19718 23704 19751
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23676 17898 23704 19450
rect 23584 17870 23704 17898
rect 23584 17338 23612 17870
rect 23664 17808 23716 17814
rect 23662 17776 23664 17785
rect 23716 17776 23718 17785
rect 23662 17711 23718 17720
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23662 17096 23718 17105
rect 23662 17031 23664 17040
rect 23716 17031 23718 17040
rect 23664 17002 23716 17008
rect 23664 16584 23716 16590
rect 23216 16561 23336 16574
rect 23202 16552 23336 16561
rect 23258 16546 23336 16552
rect 23202 16487 23258 16496
rect 23308 14958 23336 16546
rect 23664 16526 23716 16532
rect 23480 16448 23532 16454
rect 23676 16425 23704 16526
rect 23768 16522 23796 21490
rect 23860 16998 23888 23462
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 23480 16390 23532 16396
rect 23662 16416 23718 16425
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23400 15065 23428 15438
rect 23386 15056 23442 15065
rect 23386 14991 23442 15000
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22204 14278 22232 14350
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 21654 14172 21962 14181
rect 21654 14170 21660 14172
rect 21716 14170 21740 14172
rect 21796 14170 21820 14172
rect 21876 14170 21900 14172
rect 21956 14170 21962 14172
rect 21716 14118 21718 14170
rect 21898 14118 21900 14170
rect 21654 14116 21660 14118
rect 21716 14116 21740 14118
rect 21796 14116 21820 14118
rect 21876 14116 21900 14118
rect 21956 14116 21962 14118
rect 21654 14107 21962 14116
rect 20994 13628 21302 13637
rect 20994 13626 21000 13628
rect 21056 13626 21080 13628
rect 21136 13626 21160 13628
rect 21216 13626 21240 13628
rect 21296 13626 21302 13628
rect 21056 13574 21058 13626
rect 21238 13574 21240 13626
rect 20994 13572 21000 13574
rect 21056 13572 21080 13574
rect 21136 13572 21160 13574
rect 21216 13572 21240 13574
rect 21296 13572 21302 13574
rect 20994 13563 21302 13572
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19168 12986 19196 13126
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19444 12918 19472 13262
rect 19996 12918 20024 13330
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20640 12986 20668 13262
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12986 20760 13126
rect 21654 13084 21962 13093
rect 21654 13082 21660 13084
rect 21716 13082 21740 13084
rect 21796 13082 21820 13084
rect 21876 13082 21900 13084
rect 21956 13082 21962 13084
rect 21716 13030 21718 13082
rect 21898 13030 21900 13082
rect 21654 13028 21660 13030
rect 21716 13028 21740 13030
rect 21796 13028 21820 13030
rect 21876 13028 21900 13030
rect 21956 13028 21962 13030
rect 21654 13019 21962 13028
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19076 12434 19104 12718
rect 19076 12406 19196 12434
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18984 11762 19012 12242
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18524 11626 18552 11698
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 10810 18368 10950
rect 18432 10810 18460 11494
rect 18524 11354 18552 11562
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18708 10810 18736 11086
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 19168 10606 19196 12406
rect 19444 12306 19472 12854
rect 19996 12374 20024 12854
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 20916 12306 20944 12582
rect 20994 12540 21302 12549
rect 20994 12538 21000 12540
rect 21056 12538 21080 12540
rect 21136 12538 21160 12540
rect 21216 12538 21240 12540
rect 21296 12538 21302 12540
rect 21056 12486 21058 12538
rect 21238 12486 21240 12538
rect 20994 12484 21000 12486
rect 21056 12484 21080 12486
rect 21136 12484 21160 12486
rect 21216 12484 21240 12486
rect 21296 12484 21302 12486
rect 20994 12475 21302 12484
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 21376 12238 21404 12786
rect 22204 12306 22232 14214
rect 23204 13728 23256 13734
rect 23204 13670 23256 13676
rect 23216 13462 23244 13670
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 23308 13274 23336 14894
rect 23492 14414 23520 16390
rect 23662 16351 23718 16360
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23584 15026 23612 15846
rect 23676 15745 23704 16050
rect 23662 15736 23718 15745
rect 23662 15671 23718 15680
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23676 14618 23704 15302
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23662 14376 23718 14385
rect 23662 14311 23718 14320
rect 23676 13938 23704 14311
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23400 13705 23428 13874
rect 23386 13696 23442 13705
rect 23386 13631 23442 13640
rect 23216 13246 23336 13274
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23216 12714 23244 13246
rect 23676 13025 23704 13262
rect 23662 13016 23718 13025
rect 23662 12951 23718 12960
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23204 12708 23256 12714
rect 23204 12650 23256 12656
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11830 20208 12038
rect 21654 11996 21962 12005
rect 21654 11994 21660 11996
rect 21716 11994 21740 11996
rect 21796 11994 21820 11996
rect 21876 11994 21900 11996
rect 21956 11994 21962 11996
rect 21716 11942 21718 11994
rect 21898 11942 21900 11994
rect 21654 11940 21660 11942
rect 21716 11940 21740 11942
rect 21796 11940 21820 11942
rect 21876 11940 21900 11942
rect 21956 11940 21962 11942
rect 21654 11931 21962 11940
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9654 17724 9998
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17880 9722 17908 9862
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17972 9586 18000 9862
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 15927 8732 16235 8741
rect 15927 8730 15933 8732
rect 15989 8730 16013 8732
rect 16069 8730 16093 8732
rect 16149 8730 16173 8732
rect 16229 8730 16235 8732
rect 15989 8678 15991 8730
rect 16171 8678 16173 8730
rect 15927 8676 15933 8678
rect 15989 8676 16013 8678
rect 16069 8676 16093 8678
rect 16149 8676 16173 8678
rect 16229 8676 16235 8678
rect 15927 8667 16235 8676
rect 16408 8430 16436 8978
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15660 8016 15712 8022
rect 15660 7958 15712 7964
rect 16592 7954 16620 9522
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 16868 8566 16896 9318
rect 17420 8974 17448 9318
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17420 8634 17448 8910
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 16684 8090 16712 8434
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15212 7410 15240 7754
rect 15580 7410 15608 7890
rect 16684 7886 16712 8026
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 15927 7644 16235 7653
rect 15927 7642 15933 7644
rect 15989 7642 16013 7644
rect 16069 7642 16093 7644
rect 16149 7642 16173 7644
rect 16229 7642 16235 7644
rect 15989 7590 15991 7642
rect 16171 7590 16173 7642
rect 15927 7588 15933 7590
rect 15989 7588 16013 7590
rect 16069 7588 16093 7590
rect 16149 7588 16173 7590
rect 16229 7588 16235 7590
rect 15927 7579 16235 7588
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 15212 7154 15240 7346
rect 15120 7126 15240 7154
rect 15120 7018 15148 7126
rect 15267 7100 15575 7109
rect 15267 7098 15273 7100
rect 15329 7098 15353 7100
rect 15409 7098 15433 7100
rect 15489 7098 15513 7100
rect 15569 7098 15575 7100
rect 15329 7046 15331 7098
rect 15511 7046 15513 7098
rect 15267 7044 15273 7046
rect 15329 7044 15353 7046
rect 15409 7044 15433 7046
rect 15489 7044 15513 7046
rect 15569 7044 15575 7046
rect 15267 7035 15575 7044
rect 15120 6990 15240 7018
rect 16316 7002 16344 7346
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 15212 6662 15240 6990
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 6458 15516 6598
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15267 6012 15575 6021
rect 15267 6010 15273 6012
rect 15329 6010 15353 6012
rect 15409 6010 15433 6012
rect 15489 6010 15513 6012
rect 15569 6010 15575 6012
rect 15329 5958 15331 6010
rect 15511 5958 15513 6010
rect 15267 5956 15273 5958
rect 15329 5956 15353 5958
rect 15409 5956 15433 5958
rect 15489 5956 15513 5958
rect 15569 5956 15575 5958
rect 15267 5947 15575 5956
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14752 3738 14780 5170
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14844 4622 14872 5102
rect 15267 4924 15575 4933
rect 15267 4922 15273 4924
rect 15329 4922 15353 4924
rect 15409 4922 15433 4924
rect 15489 4922 15513 4924
rect 15569 4922 15575 4924
rect 15329 4870 15331 4922
rect 15511 4870 15513 4922
rect 15267 4868 15273 4870
rect 15329 4868 15353 4870
rect 15409 4868 15433 4870
rect 15489 4868 15513 4870
rect 15569 4868 15575 4870
rect 15267 4859 15575 4868
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14844 4078 14872 4558
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 15108 4072 15160 4078
rect 15672 4026 15700 6666
rect 15927 6556 16235 6565
rect 15927 6554 15933 6556
rect 15989 6554 16013 6556
rect 16069 6554 16093 6556
rect 16149 6554 16173 6556
rect 16229 6554 16235 6556
rect 15989 6502 15991 6554
rect 16171 6502 16173 6554
rect 15927 6500 15933 6502
rect 15989 6500 16013 6502
rect 16069 6500 16093 6502
rect 16149 6500 16173 6502
rect 16229 6500 16235 6502
rect 15927 6491 16235 6500
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15764 5166 15792 6258
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15764 4758 15792 4966
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 15856 4162 15884 6054
rect 15927 5468 16235 5477
rect 15927 5466 15933 5468
rect 15989 5466 16013 5468
rect 16069 5466 16093 5468
rect 16149 5466 16173 5468
rect 16229 5466 16235 5468
rect 15989 5414 15991 5466
rect 16171 5414 16173 5466
rect 15927 5412 15933 5414
rect 15989 5412 16013 5414
rect 16069 5412 16093 5414
rect 16149 5412 16173 5414
rect 16229 5412 16235 5414
rect 15927 5403 16235 5412
rect 15927 4380 16235 4389
rect 15927 4378 15933 4380
rect 15989 4378 16013 4380
rect 16069 4378 16093 4380
rect 16149 4378 16173 4380
rect 16229 4378 16235 4380
rect 15989 4326 15991 4378
rect 16171 4326 16173 4378
rect 15927 4324 15933 4326
rect 15989 4324 16013 4326
rect 16069 4324 16093 4326
rect 16149 4324 16173 4326
rect 16229 4324 16235 4326
rect 15927 4315 16235 4324
rect 15108 4014 15160 4020
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14844 3602 14872 3878
rect 15120 3754 15148 4014
rect 15580 4010 15700 4026
rect 15568 4004 15700 4010
rect 15620 3998 15700 4004
rect 15764 4134 15884 4162
rect 15568 3946 15620 3952
rect 15267 3836 15575 3845
rect 15267 3834 15273 3836
rect 15329 3834 15353 3836
rect 15409 3834 15433 3836
rect 15489 3834 15513 3836
rect 15569 3834 15575 3836
rect 15329 3782 15331 3834
rect 15511 3782 15513 3834
rect 15267 3780 15273 3782
rect 15329 3780 15353 3782
rect 15409 3780 15433 3782
rect 15489 3780 15513 3782
rect 15569 3780 15575 3782
rect 15267 3771 15575 3780
rect 15120 3738 15240 3754
rect 15120 3732 15252 3738
rect 15120 3726 15200 3732
rect 15200 3674 15252 3680
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14844 3466 14872 3538
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 3194 14872 3402
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15028 2854 15056 2994
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 15028 2446 15056 2790
rect 15120 2650 15148 2926
rect 15267 2748 15575 2757
rect 15267 2746 15273 2748
rect 15329 2746 15353 2748
rect 15409 2746 15433 2748
rect 15489 2746 15513 2748
rect 15569 2746 15575 2748
rect 15329 2694 15331 2746
rect 15511 2694 15513 2746
rect 15267 2692 15273 2694
rect 15329 2692 15353 2694
rect 15409 2692 15433 2694
rect 15489 2692 15513 2694
rect 15569 2692 15575 2694
rect 15267 2683 15575 2692
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 15568 2440 15620 2446
rect 15672 2428 15700 2994
rect 15764 2774 15792 4134
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15856 3534 15884 4014
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15856 3194 15884 3470
rect 15927 3292 16235 3301
rect 15927 3290 15933 3292
rect 15989 3290 16013 3292
rect 16069 3290 16093 3292
rect 16149 3290 16173 3292
rect 16229 3290 16235 3292
rect 15989 3238 15991 3290
rect 16171 3238 16173 3290
rect 15927 3236 15933 3238
rect 15989 3236 16013 3238
rect 16069 3236 16093 3238
rect 16149 3236 16173 3238
rect 16229 3236 16235 3238
rect 15927 3227 16235 3236
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15764 2746 15884 2774
rect 15856 2446 15884 2746
rect 15948 2650 15976 2926
rect 16040 2650 16068 3062
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16408 2446 16436 7210
rect 16500 2582 16528 7686
rect 16960 6866 16988 7890
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 4010 16712 6598
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 17052 2446 17080 7142
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 5914 17264 6598
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17604 5710 17632 6054
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17604 5250 17632 5646
rect 17512 5222 17632 5250
rect 17868 5228 17920 5234
rect 17512 5166 17540 5222
rect 17868 5170 17920 5176
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17604 3738 17632 4082
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17696 3738 17724 4014
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17880 3602 17908 5170
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17512 2582 17540 2790
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 17972 2446 18000 8298
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 18156 6254 18184 6870
rect 18248 6458 18276 8434
rect 18524 8430 18552 10066
rect 19168 9874 19196 10542
rect 19260 10130 19288 11154
rect 20732 10674 20760 11494
rect 20994 11452 21302 11461
rect 20994 11450 21000 11452
rect 21056 11450 21080 11452
rect 21136 11450 21160 11452
rect 21216 11450 21240 11452
rect 21296 11450 21302 11452
rect 21056 11398 21058 11450
rect 21238 11398 21240 11450
rect 20994 11396 21000 11398
rect 21056 11396 21080 11398
rect 21136 11396 21160 11398
rect 21216 11396 21240 11398
rect 21296 11396 21302 11398
rect 20994 11387 21302 11396
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 19616 10532 19668 10538
rect 19616 10474 19668 10480
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19628 10062 19656 10474
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 19996 10130 20024 10406
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19352 9874 19380 9930
rect 19168 9846 19380 9874
rect 19260 9042 19288 9846
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18708 6866 18736 7346
rect 19076 7342 19104 8434
rect 19260 8430 19288 8978
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18892 6798 18920 7278
rect 19260 6934 19288 8366
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18524 6390 18552 6598
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18064 5166 18092 5714
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18064 4078 18092 5102
rect 18156 4282 18184 6190
rect 18892 6186 18920 6734
rect 19260 6390 19288 6870
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18984 5846 19012 6258
rect 19168 5914 19196 6258
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19260 5914 19288 6190
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 19996 5710 20024 6258
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19996 5370 20024 5646
rect 20180 5642 20208 6190
rect 20168 5636 20220 5642
rect 20168 5578 20220 5584
rect 20180 5370 20208 5578
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18156 3670 18184 4082
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18340 3738 18368 4014
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18156 3466 18184 3606
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 18156 3194 18184 3402
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18248 2990 18276 3402
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 3194 18828 3334
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 19536 3058 19564 3402
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 2650 19472 2926
rect 19536 2650 19564 2994
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 20272 2446 20300 10134
rect 20456 10062 20484 10406
rect 20732 10130 20760 10610
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20916 10266 20944 10542
rect 20994 10364 21302 10373
rect 20994 10362 21000 10364
rect 21056 10362 21080 10364
rect 21136 10362 21160 10364
rect 21216 10362 21240 10364
rect 21296 10362 21302 10364
rect 21056 10310 21058 10362
rect 21238 10310 21240 10362
rect 20994 10308 21000 10310
rect 21056 10308 21080 10310
rect 21136 10308 21160 10310
rect 21216 10308 21240 10310
rect 21296 10308 21302 10310
rect 20994 10299 21302 10308
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20994 9276 21302 9285
rect 20994 9274 21000 9276
rect 21056 9274 21080 9276
rect 21136 9274 21160 9276
rect 21216 9274 21240 9276
rect 21296 9274 21302 9276
rect 21056 9222 21058 9274
rect 21238 9222 21240 9274
rect 20994 9220 21000 9222
rect 21056 9220 21080 9222
rect 21136 9220 21160 9222
rect 21216 9220 21240 9222
rect 21296 9220 21302 9222
rect 20994 9211 21302 9220
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20364 4826 20392 5102
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20456 2922 20484 5102
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20732 2774 20760 8298
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20916 7954 20944 8230
rect 20994 8188 21302 8197
rect 20994 8186 21000 8188
rect 21056 8186 21080 8188
rect 21136 8186 21160 8188
rect 21216 8186 21240 8188
rect 21296 8186 21302 8188
rect 21056 8134 21058 8186
rect 21238 8134 21240 8186
rect 20994 8132 21000 8134
rect 21056 8132 21080 8134
rect 21136 8132 21160 8134
rect 21216 8132 21240 8134
rect 21296 8132 21302 8134
rect 20994 8123 21302 8132
rect 21376 8022 21404 11018
rect 21468 10266 21496 11018
rect 21560 10606 21588 11086
rect 21654 10908 21962 10917
rect 21654 10906 21660 10908
rect 21716 10906 21740 10908
rect 21796 10906 21820 10908
rect 21876 10906 21900 10908
rect 21956 10906 21962 10908
rect 21716 10854 21718 10906
rect 21898 10854 21900 10906
rect 21654 10852 21660 10854
rect 21716 10852 21740 10854
rect 21796 10852 21820 10854
rect 21876 10852 21900 10854
rect 21956 10852 21962 10854
rect 21654 10843 21962 10852
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21560 9994 21588 10542
rect 21652 10062 21680 10610
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10266 22048 10542
rect 22112 10266 22140 10610
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22204 10198 22232 12242
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22664 10470 22692 11154
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22664 10130 22692 10406
rect 23032 10130 23060 10950
rect 23216 10606 23244 12650
rect 23400 12345 23428 12786
rect 23386 12336 23442 12345
rect 23386 12271 23442 12280
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23676 11665 23704 11698
rect 23662 11656 23718 11665
rect 23662 11591 23718 11600
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21654 9820 21962 9829
rect 21654 9818 21660 9820
rect 21716 9818 21740 9820
rect 21796 9818 21820 9820
rect 21876 9818 21900 9820
rect 21956 9818 21962 9820
rect 21716 9766 21718 9818
rect 21898 9766 21900 9818
rect 21654 9764 21660 9766
rect 21716 9764 21740 9766
rect 21796 9764 21820 9766
rect 21876 9764 21900 9766
rect 21956 9764 21962 9766
rect 21654 9755 21962 9764
rect 21654 8732 21962 8741
rect 21654 8730 21660 8732
rect 21716 8730 21740 8732
rect 21796 8730 21820 8732
rect 21876 8730 21900 8732
rect 21956 8730 21962 8732
rect 21716 8678 21718 8730
rect 21898 8678 21900 8730
rect 21654 8676 21660 8678
rect 21716 8676 21740 8678
rect 21796 8676 21820 8678
rect 21876 8676 21900 8678
rect 21956 8676 21962 8678
rect 21654 8667 21962 8676
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 7342 21128 7686
rect 21376 7410 21404 7958
rect 21744 7954 21772 8230
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21548 7812 21600 7818
rect 21548 7754 21600 7760
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 20994 7100 21302 7109
rect 20994 7098 21000 7100
rect 21056 7098 21080 7100
rect 21136 7098 21160 7100
rect 21216 7098 21240 7100
rect 21296 7098 21302 7100
rect 21056 7046 21058 7098
rect 21238 7046 21240 7098
rect 20994 7044 21000 7046
rect 21056 7044 21080 7046
rect 21136 7044 21160 7046
rect 21216 7044 21240 7046
rect 21296 7044 21302 7046
rect 20994 7035 21302 7044
rect 21560 6934 21588 7754
rect 21654 7644 21962 7653
rect 21654 7642 21660 7644
rect 21716 7642 21740 7644
rect 21796 7642 21820 7644
rect 21876 7642 21900 7644
rect 21956 7642 21962 7644
rect 21716 7590 21718 7642
rect 21898 7590 21900 7642
rect 21654 7588 21660 7590
rect 21716 7588 21740 7590
rect 21796 7588 21820 7590
rect 21876 7588 21900 7590
rect 21956 7588 21962 7590
rect 21654 7579 21962 7588
rect 22020 7342 22048 7754
rect 22112 7342 22140 8026
rect 22204 7886 22232 8230
rect 22480 8090 22508 8366
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 20994 6012 21302 6021
rect 20994 6010 21000 6012
rect 21056 6010 21080 6012
rect 21136 6010 21160 6012
rect 21216 6010 21240 6012
rect 21296 6010 21302 6012
rect 21056 5958 21058 6010
rect 21238 5958 21240 6010
rect 20994 5956 21000 5958
rect 21056 5956 21080 5958
rect 21136 5956 21160 5958
rect 21216 5956 21240 5958
rect 21296 5956 21302 5958
rect 20994 5947 21302 5956
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 20824 4706 20852 5170
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20916 4826 20944 5102
rect 20994 4924 21302 4933
rect 20994 4922 21000 4924
rect 21056 4922 21080 4924
rect 21136 4922 21160 4924
rect 21216 4922 21240 4924
rect 21296 4922 21302 4924
rect 21056 4870 21058 4922
rect 21238 4870 21240 4922
rect 20994 4868 21000 4870
rect 21056 4868 21080 4870
rect 21136 4868 21160 4870
rect 21216 4868 21240 4870
rect 21296 4868 21302 4870
rect 20994 4859 21302 4868
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20824 4678 20944 4706
rect 20916 4554 20944 4678
rect 21376 4622 21404 5170
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 20916 3738 20944 4490
rect 20994 3836 21302 3845
rect 20994 3834 21000 3836
rect 21056 3834 21080 3836
rect 21136 3834 21160 3836
rect 21216 3834 21240 3836
rect 21296 3834 21302 3836
rect 21056 3782 21058 3834
rect 21238 3782 21240 3834
rect 20994 3780 21000 3782
rect 21056 3780 21080 3782
rect 21136 3780 21160 3782
rect 21216 3780 21240 3782
rect 21296 3780 21302 3782
rect 20994 3771 21302 3780
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 21468 3602 21496 5102
rect 21560 4690 21588 6870
rect 22112 6866 22140 7278
rect 22204 6934 22232 7346
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22480 6798 22508 7686
rect 22572 7546 22600 8434
rect 22940 7546 22968 8434
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 7546 23060 8230
rect 23124 7954 23152 10066
rect 23112 7948 23164 7954
rect 23112 7890 23164 7896
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 21654 6556 21962 6565
rect 21654 6554 21660 6556
rect 21716 6554 21740 6556
rect 21796 6554 21820 6556
rect 21876 6554 21900 6556
rect 21956 6554 21962 6556
rect 21716 6502 21718 6554
rect 21898 6502 21900 6554
rect 21654 6500 21660 6502
rect 21716 6500 21740 6502
rect 21796 6500 21820 6502
rect 21876 6500 21900 6502
rect 21956 6500 21962 6502
rect 21654 6491 21962 6500
rect 21654 5468 21962 5477
rect 21654 5466 21660 5468
rect 21716 5466 21740 5468
rect 21796 5466 21820 5468
rect 21876 5466 21900 5468
rect 21956 5466 21962 5468
rect 21716 5414 21718 5466
rect 21898 5414 21900 5466
rect 21654 5412 21660 5414
rect 21716 5412 21740 5414
rect 21796 5412 21820 5414
rect 21876 5412 21900 5414
rect 21956 5412 21962 5414
rect 21654 5403 21962 5412
rect 23124 5166 23152 7890
rect 23216 7342 23244 10542
rect 23308 9926 23336 11086
rect 23400 10985 23428 11086
rect 23386 10976 23442 10985
rect 23386 10911 23442 10920
rect 23662 10296 23718 10305
rect 23662 10231 23718 10240
rect 23676 10062 23704 10231
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23308 5914 23336 9862
rect 23572 9716 23624 9722
rect 23572 9658 23624 9664
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23400 8265 23428 8298
rect 23386 8256 23442 8265
rect 23386 8191 23442 8200
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23492 6458 23520 7822
rect 23584 6798 23612 9658
rect 23662 9616 23718 9625
rect 23662 9551 23718 9560
rect 23676 9450 23704 9551
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23662 8936 23718 8945
rect 23662 8871 23718 8880
rect 23676 8838 23704 8871
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23662 7576 23718 7585
rect 23662 7511 23718 7520
rect 23676 7410 23704 7511
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23662 6896 23718 6905
rect 23662 6831 23718 6840
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23676 6662 23704 6831
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23676 6225 23704 6258
rect 23662 6216 23718 6225
rect 23662 6151 23718 6160
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23400 5545 23428 5646
rect 23386 5536 23442 5545
rect 23386 5471 23442 5480
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 23112 5160 23164 5166
rect 23112 5102 23164 5108
rect 23676 4865 23704 5170
rect 23662 4856 23718 4865
rect 23662 4791 23718 4800
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23664 4616 23716 4622
rect 23664 4558 23716 4564
rect 21654 4380 21962 4389
rect 21654 4378 21660 4380
rect 21716 4378 21740 4380
rect 21796 4378 21820 4380
rect 21876 4378 21900 4380
rect 21956 4378 21962 4380
rect 21716 4326 21718 4378
rect 21898 4326 21900 4378
rect 21654 4324 21660 4326
rect 21716 4324 21740 4326
rect 21796 4324 21820 4326
rect 21876 4324 21900 4326
rect 21956 4324 21962 4326
rect 21654 4315 21962 4324
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21654 3292 21962 3301
rect 21654 3290 21660 3292
rect 21716 3290 21740 3292
rect 21796 3290 21820 3292
rect 21876 3290 21900 3292
rect 21956 3290 21962 3292
rect 21716 3238 21718 3290
rect 21898 3238 21900 3290
rect 21654 3236 21660 3238
rect 21716 3236 21740 3238
rect 21796 3236 21820 3238
rect 21876 3236 21900 3238
rect 21956 3236 21962 3238
rect 21654 3227 21962 3236
rect 23492 3194 23520 4558
rect 23676 4185 23704 4558
rect 23662 4176 23718 4185
rect 23662 4111 23718 4120
rect 23664 3528 23716 3534
rect 23662 3496 23664 3505
rect 23716 3496 23718 3505
rect 23662 3431 23718 3440
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23676 2825 23704 2994
rect 23662 2816 23718 2825
rect 20732 2746 20852 2774
rect 20824 2446 20852 2746
rect 20994 2748 21302 2757
rect 23662 2751 23718 2760
rect 20994 2746 21000 2748
rect 21056 2746 21080 2748
rect 21136 2746 21160 2748
rect 21216 2746 21240 2748
rect 21296 2746 21302 2748
rect 21056 2694 21058 2746
rect 21238 2694 21240 2746
rect 20994 2692 21000 2694
rect 21056 2692 21080 2694
rect 21136 2692 21160 2694
rect 21216 2692 21240 2694
rect 21296 2692 21302 2694
rect 20994 2683 21302 2692
rect 15620 2400 15700 2428
rect 15844 2440 15896 2446
rect 15568 2382 15620 2388
rect 15844 2382 15896 2388
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 10980 800 11008 2382
rect 11624 800 11652 2382
rect 12268 800 12296 2382
rect 12912 800 12940 2382
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 800 13584 2246
rect 14200 800 14228 2382
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 14844 800 14872 2314
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 15580 1170 15608 2246
rect 15927 2204 16235 2213
rect 15927 2202 15933 2204
rect 15989 2202 16013 2204
rect 16069 2202 16093 2204
rect 16149 2202 16173 2204
rect 16229 2202 16235 2204
rect 15989 2150 15991 2202
rect 16171 2150 16173 2202
rect 15927 2148 15933 2150
rect 15989 2148 16013 2150
rect 16069 2148 16093 2150
rect 16149 2148 16173 2150
rect 16229 2148 16235 2150
rect 15927 2139 16235 2148
rect 16316 1170 16344 2246
rect 15488 1142 15608 1170
rect 16132 1142 16344 1170
rect 15488 800 15516 1142
rect 16132 800 16160 1142
rect 16776 800 16804 2246
rect 17420 800 17448 2382
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 800 18092 2246
rect 18708 800 18736 2382
rect 19352 800 19380 2382
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 19996 800 20024 2246
rect 20640 800 20668 2246
rect 21284 800 21312 2382
rect 21654 2204 21962 2213
rect 21654 2202 21660 2204
rect 21716 2202 21740 2204
rect 21796 2202 21820 2204
rect 21876 2202 21900 2204
rect 21956 2202 21962 2204
rect 21716 2150 21718 2202
rect 21898 2150 21900 2202
rect 21654 2148 21660 2150
rect 21716 2148 21740 2150
rect 21796 2148 21820 2150
rect 21876 2148 21900 2150
rect 21956 2148 21962 2150
rect 21654 2139 21962 2148
rect 10428 734 10640 762
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
<< via2 >>
rect 4479 25050 4535 25052
rect 4559 25050 4615 25052
rect 4639 25050 4695 25052
rect 4719 25050 4775 25052
rect 4479 24998 4525 25050
rect 4525 24998 4535 25050
rect 4559 24998 4589 25050
rect 4589 24998 4601 25050
rect 4601 24998 4615 25050
rect 4639 24998 4653 25050
rect 4653 24998 4665 25050
rect 4665 24998 4695 25050
rect 4719 24998 4729 25050
rect 4729 24998 4775 25050
rect 4479 24996 4535 24998
rect 4559 24996 4615 24998
rect 4639 24996 4695 24998
rect 4719 24996 4775 24998
rect 3819 24506 3875 24508
rect 3899 24506 3955 24508
rect 3979 24506 4035 24508
rect 4059 24506 4115 24508
rect 3819 24454 3865 24506
rect 3865 24454 3875 24506
rect 3899 24454 3929 24506
rect 3929 24454 3941 24506
rect 3941 24454 3955 24506
rect 3979 24454 3993 24506
rect 3993 24454 4005 24506
rect 4005 24454 4035 24506
rect 4059 24454 4069 24506
rect 4069 24454 4115 24506
rect 3819 24452 3875 24454
rect 3899 24452 3955 24454
rect 3979 24452 4035 24454
rect 4059 24452 4115 24454
rect 4479 23962 4535 23964
rect 4559 23962 4615 23964
rect 4639 23962 4695 23964
rect 4719 23962 4775 23964
rect 4479 23910 4525 23962
rect 4525 23910 4535 23962
rect 4559 23910 4589 23962
rect 4589 23910 4601 23962
rect 4601 23910 4615 23962
rect 4639 23910 4653 23962
rect 4653 23910 4665 23962
rect 4665 23910 4695 23962
rect 4719 23910 4729 23962
rect 4729 23910 4775 23962
rect 4479 23908 4535 23910
rect 4559 23908 4615 23910
rect 4639 23908 4695 23910
rect 4719 23908 4775 23910
rect 3819 23418 3875 23420
rect 3899 23418 3955 23420
rect 3979 23418 4035 23420
rect 4059 23418 4115 23420
rect 3819 23366 3865 23418
rect 3865 23366 3875 23418
rect 3899 23366 3929 23418
rect 3929 23366 3941 23418
rect 3941 23366 3955 23418
rect 3979 23366 3993 23418
rect 3993 23366 4005 23418
rect 4005 23366 4035 23418
rect 4059 23366 4069 23418
rect 4069 23366 4115 23418
rect 3819 23364 3875 23366
rect 3899 23364 3955 23366
rect 3979 23364 4035 23366
rect 4059 23364 4115 23366
rect 4479 22874 4535 22876
rect 4559 22874 4615 22876
rect 4639 22874 4695 22876
rect 4719 22874 4775 22876
rect 4479 22822 4525 22874
rect 4525 22822 4535 22874
rect 4559 22822 4589 22874
rect 4589 22822 4601 22874
rect 4601 22822 4615 22874
rect 4639 22822 4653 22874
rect 4653 22822 4665 22874
rect 4665 22822 4695 22874
rect 4719 22822 4729 22874
rect 4729 22822 4775 22874
rect 4479 22820 4535 22822
rect 4559 22820 4615 22822
rect 4639 22820 4695 22822
rect 4719 22820 4775 22822
rect 3819 22330 3875 22332
rect 3899 22330 3955 22332
rect 3979 22330 4035 22332
rect 4059 22330 4115 22332
rect 3819 22278 3865 22330
rect 3865 22278 3875 22330
rect 3899 22278 3929 22330
rect 3929 22278 3941 22330
rect 3941 22278 3955 22330
rect 3979 22278 3993 22330
rect 3993 22278 4005 22330
rect 4005 22278 4035 22330
rect 4059 22278 4069 22330
rect 4069 22278 4115 22330
rect 3819 22276 3875 22278
rect 3899 22276 3955 22278
rect 3979 22276 4035 22278
rect 4059 22276 4115 22278
rect 4479 21786 4535 21788
rect 4559 21786 4615 21788
rect 4639 21786 4695 21788
rect 4719 21786 4775 21788
rect 4479 21734 4525 21786
rect 4525 21734 4535 21786
rect 4559 21734 4589 21786
rect 4589 21734 4601 21786
rect 4601 21734 4615 21786
rect 4639 21734 4653 21786
rect 4653 21734 4665 21786
rect 4665 21734 4695 21786
rect 4719 21734 4729 21786
rect 4729 21734 4775 21786
rect 4479 21732 4535 21734
rect 4559 21732 4615 21734
rect 4639 21732 4695 21734
rect 4719 21732 4775 21734
rect 846 21256 902 21312
rect 3819 21242 3875 21244
rect 3899 21242 3955 21244
rect 3979 21242 4035 21244
rect 4059 21242 4115 21244
rect 3819 21190 3865 21242
rect 3865 21190 3875 21242
rect 3899 21190 3929 21242
rect 3929 21190 3941 21242
rect 3941 21190 3955 21242
rect 3979 21190 3993 21242
rect 3993 21190 4005 21242
rect 4005 21190 4035 21242
rect 4059 21190 4069 21242
rect 4069 21190 4115 21242
rect 3819 21188 3875 21190
rect 3899 21188 3955 21190
rect 3979 21188 4035 21190
rect 4059 21188 4115 21190
rect 1398 20440 1454 20496
rect 846 19896 902 19952
rect 4479 20698 4535 20700
rect 4559 20698 4615 20700
rect 4639 20698 4695 20700
rect 4719 20698 4775 20700
rect 4479 20646 4525 20698
rect 4525 20646 4535 20698
rect 4559 20646 4589 20698
rect 4589 20646 4601 20698
rect 4601 20646 4615 20698
rect 4639 20646 4653 20698
rect 4653 20646 4665 20698
rect 4665 20646 4695 20698
rect 4719 20646 4729 20698
rect 4729 20646 4775 20698
rect 4479 20644 4535 20646
rect 4559 20644 4615 20646
rect 4639 20644 4695 20646
rect 4719 20644 4775 20646
rect 3819 20154 3875 20156
rect 3899 20154 3955 20156
rect 3979 20154 4035 20156
rect 4059 20154 4115 20156
rect 3819 20102 3865 20154
rect 3865 20102 3875 20154
rect 3899 20102 3929 20154
rect 3929 20102 3941 20154
rect 3941 20102 3955 20154
rect 3979 20102 3993 20154
rect 3993 20102 4005 20154
rect 4005 20102 4035 20154
rect 4059 20102 4069 20154
rect 4069 20102 4115 20154
rect 3819 20100 3875 20102
rect 3899 20100 3955 20102
rect 3979 20100 4035 20102
rect 4059 20100 4115 20102
rect 1398 19116 1400 19136
rect 1400 19116 1452 19136
rect 1452 19116 1454 19136
rect 1398 19080 1454 19116
rect 3819 19066 3875 19068
rect 3899 19066 3955 19068
rect 3979 19066 4035 19068
rect 4059 19066 4115 19068
rect 3819 19014 3865 19066
rect 3865 19014 3875 19066
rect 3899 19014 3929 19066
rect 3929 19014 3941 19066
rect 3941 19014 3955 19066
rect 3979 19014 3993 19066
rect 3993 19014 4005 19066
rect 4005 19014 4035 19066
rect 4059 19014 4069 19066
rect 4069 19014 4115 19066
rect 3819 19012 3875 19014
rect 3899 19012 3955 19014
rect 3979 19012 4035 19014
rect 4059 19012 4115 19014
rect 4479 19610 4535 19612
rect 4559 19610 4615 19612
rect 4639 19610 4695 19612
rect 4719 19610 4775 19612
rect 4479 19558 4525 19610
rect 4525 19558 4535 19610
rect 4559 19558 4589 19610
rect 4589 19558 4601 19610
rect 4601 19558 4615 19610
rect 4639 19558 4653 19610
rect 4653 19558 4665 19610
rect 4665 19558 4695 19610
rect 4719 19558 4729 19610
rect 4729 19558 4775 19610
rect 4479 19556 4535 19558
rect 4559 19556 4615 19558
rect 4639 19556 4695 19558
rect 4719 19556 4775 19558
rect 846 18572 848 18592
rect 848 18572 900 18592
rect 900 18572 902 18592
rect 846 18536 902 18572
rect 4479 18522 4535 18524
rect 4559 18522 4615 18524
rect 4639 18522 4695 18524
rect 4719 18522 4775 18524
rect 4479 18470 4525 18522
rect 4525 18470 4535 18522
rect 4559 18470 4589 18522
rect 4589 18470 4601 18522
rect 4601 18470 4615 18522
rect 4639 18470 4653 18522
rect 4653 18470 4665 18522
rect 4665 18470 4695 18522
rect 4719 18470 4729 18522
rect 4729 18470 4775 18522
rect 4479 18468 4535 18470
rect 4559 18468 4615 18470
rect 4639 18468 4695 18470
rect 4719 18468 4775 18470
rect 3819 17978 3875 17980
rect 3899 17978 3955 17980
rect 3979 17978 4035 17980
rect 4059 17978 4115 17980
rect 3819 17926 3865 17978
rect 3865 17926 3875 17978
rect 3899 17926 3929 17978
rect 3929 17926 3941 17978
rect 3941 17926 3955 17978
rect 3979 17926 3993 17978
rect 3993 17926 4005 17978
rect 4005 17926 4035 17978
rect 4059 17926 4069 17978
rect 4069 17926 4115 17978
rect 3819 17924 3875 17926
rect 3899 17924 3955 17926
rect 3979 17924 4035 17926
rect 4059 17924 4115 17926
rect 1398 17720 1454 17776
rect 846 17196 902 17232
rect 846 17176 848 17196
rect 848 17176 900 17196
rect 900 17176 902 17196
rect 3819 16890 3875 16892
rect 3899 16890 3955 16892
rect 3979 16890 4035 16892
rect 4059 16890 4115 16892
rect 3819 16838 3865 16890
rect 3865 16838 3875 16890
rect 3899 16838 3929 16890
rect 3929 16838 3941 16890
rect 3941 16838 3955 16890
rect 3979 16838 3993 16890
rect 3993 16838 4005 16890
rect 4005 16838 4035 16890
rect 4059 16838 4069 16890
rect 4069 16838 4115 16890
rect 3819 16836 3875 16838
rect 3899 16836 3955 16838
rect 3979 16836 4035 16838
rect 4059 16836 4115 16838
rect 846 16532 848 16552
rect 848 16532 900 16552
rect 900 16532 902 16552
rect 846 16496 902 16532
rect 4479 17434 4535 17436
rect 4559 17434 4615 17436
rect 4639 17434 4695 17436
rect 4719 17434 4775 17436
rect 4479 17382 4525 17434
rect 4525 17382 4535 17434
rect 4559 17382 4589 17434
rect 4589 17382 4601 17434
rect 4601 17382 4615 17434
rect 4639 17382 4653 17434
rect 4653 17382 4665 17434
rect 4665 17382 4695 17434
rect 4719 17382 4729 17434
rect 4729 17382 4775 17434
rect 4479 17380 4535 17382
rect 4559 17380 4615 17382
rect 4639 17380 4695 17382
rect 4719 17380 4775 17382
rect 4479 16346 4535 16348
rect 4559 16346 4615 16348
rect 4639 16346 4695 16348
rect 4719 16346 4775 16348
rect 4479 16294 4525 16346
rect 4525 16294 4535 16346
rect 4559 16294 4589 16346
rect 4589 16294 4601 16346
rect 4601 16294 4615 16346
rect 4639 16294 4653 16346
rect 4653 16294 4665 16346
rect 4665 16294 4695 16346
rect 4719 16294 4729 16346
rect 4729 16294 4775 16346
rect 4479 16292 4535 16294
rect 4559 16292 4615 16294
rect 4639 16292 4695 16294
rect 4719 16292 4775 16294
rect 846 15816 902 15872
rect 3819 15802 3875 15804
rect 3899 15802 3955 15804
rect 3979 15802 4035 15804
rect 4059 15802 4115 15804
rect 3819 15750 3865 15802
rect 3865 15750 3875 15802
rect 3899 15750 3929 15802
rect 3929 15750 3941 15802
rect 3941 15750 3955 15802
rect 3979 15750 3993 15802
rect 3993 15750 4005 15802
rect 4005 15750 4035 15802
rect 4059 15750 4069 15802
rect 4069 15750 4115 15802
rect 3819 15748 3875 15750
rect 3899 15748 3955 15750
rect 3979 15748 4035 15750
rect 4059 15748 4115 15750
rect 10206 25050 10262 25052
rect 10286 25050 10342 25052
rect 10366 25050 10422 25052
rect 10446 25050 10502 25052
rect 10206 24998 10252 25050
rect 10252 24998 10262 25050
rect 10286 24998 10316 25050
rect 10316 24998 10328 25050
rect 10328 24998 10342 25050
rect 10366 24998 10380 25050
rect 10380 24998 10392 25050
rect 10392 24998 10422 25050
rect 10446 24998 10456 25050
rect 10456 24998 10502 25050
rect 10206 24996 10262 24998
rect 10286 24996 10342 24998
rect 10366 24996 10422 24998
rect 10446 24996 10502 24998
rect 9546 24506 9602 24508
rect 9626 24506 9682 24508
rect 9706 24506 9762 24508
rect 9786 24506 9842 24508
rect 9546 24454 9592 24506
rect 9592 24454 9602 24506
rect 9626 24454 9656 24506
rect 9656 24454 9668 24506
rect 9668 24454 9682 24506
rect 9706 24454 9720 24506
rect 9720 24454 9732 24506
rect 9732 24454 9762 24506
rect 9786 24454 9796 24506
rect 9796 24454 9842 24506
rect 9546 24452 9602 24454
rect 9626 24452 9682 24454
rect 9706 24452 9762 24454
rect 9786 24452 9842 24454
rect 9546 23418 9602 23420
rect 9626 23418 9682 23420
rect 9706 23418 9762 23420
rect 9786 23418 9842 23420
rect 9546 23366 9592 23418
rect 9592 23366 9602 23418
rect 9626 23366 9656 23418
rect 9656 23366 9668 23418
rect 9668 23366 9682 23418
rect 9706 23366 9720 23418
rect 9720 23366 9732 23418
rect 9732 23366 9762 23418
rect 9786 23366 9796 23418
rect 9796 23366 9842 23418
rect 9546 23364 9602 23366
rect 9626 23364 9682 23366
rect 9706 23364 9762 23366
rect 9786 23364 9842 23366
rect 9546 22330 9602 22332
rect 9626 22330 9682 22332
rect 9706 22330 9762 22332
rect 9786 22330 9842 22332
rect 9546 22278 9592 22330
rect 9592 22278 9602 22330
rect 9626 22278 9656 22330
rect 9656 22278 9668 22330
rect 9668 22278 9682 22330
rect 9706 22278 9720 22330
rect 9720 22278 9732 22330
rect 9732 22278 9762 22330
rect 9786 22278 9796 22330
rect 9796 22278 9842 22330
rect 9546 22276 9602 22278
rect 9626 22276 9682 22278
rect 9706 22276 9762 22278
rect 9786 22276 9842 22278
rect 9546 21242 9602 21244
rect 9626 21242 9682 21244
rect 9706 21242 9762 21244
rect 9786 21242 9842 21244
rect 9546 21190 9592 21242
rect 9592 21190 9602 21242
rect 9626 21190 9656 21242
rect 9656 21190 9668 21242
rect 9668 21190 9682 21242
rect 9706 21190 9720 21242
rect 9720 21190 9732 21242
rect 9732 21190 9762 21242
rect 9786 21190 9796 21242
rect 9796 21190 9842 21242
rect 9546 21188 9602 21190
rect 9626 21188 9682 21190
rect 9706 21188 9762 21190
rect 9786 21188 9842 21190
rect 9546 20154 9602 20156
rect 9626 20154 9682 20156
rect 9706 20154 9762 20156
rect 9786 20154 9842 20156
rect 9546 20102 9592 20154
rect 9592 20102 9602 20154
rect 9626 20102 9656 20154
rect 9656 20102 9668 20154
rect 9668 20102 9682 20154
rect 9706 20102 9720 20154
rect 9720 20102 9732 20154
rect 9732 20102 9762 20154
rect 9786 20102 9796 20154
rect 9796 20102 9842 20154
rect 9546 20100 9602 20102
rect 9626 20100 9682 20102
rect 9706 20100 9762 20102
rect 9786 20100 9842 20102
rect 9546 19066 9602 19068
rect 9626 19066 9682 19068
rect 9706 19066 9762 19068
rect 9786 19066 9842 19068
rect 9546 19014 9592 19066
rect 9592 19014 9602 19066
rect 9626 19014 9656 19066
rect 9656 19014 9668 19066
rect 9668 19014 9682 19066
rect 9706 19014 9720 19066
rect 9720 19014 9732 19066
rect 9732 19014 9762 19066
rect 9786 19014 9796 19066
rect 9796 19014 9842 19066
rect 9546 19012 9602 19014
rect 9626 19012 9682 19014
rect 9706 19012 9762 19014
rect 9786 19012 9842 19014
rect 1398 15000 1454 15056
rect 4479 15258 4535 15260
rect 4559 15258 4615 15260
rect 4639 15258 4695 15260
rect 4719 15258 4775 15260
rect 4479 15206 4525 15258
rect 4525 15206 4535 15258
rect 4559 15206 4589 15258
rect 4589 15206 4601 15258
rect 4601 15206 4615 15258
rect 4639 15206 4653 15258
rect 4653 15206 4665 15258
rect 4665 15206 4695 15258
rect 4719 15206 4729 15258
rect 4729 15206 4775 15258
rect 4479 15204 4535 15206
rect 4559 15204 4615 15206
rect 4639 15204 4695 15206
rect 4719 15204 4775 15206
rect 3819 14714 3875 14716
rect 3899 14714 3955 14716
rect 3979 14714 4035 14716
rect 4059 14714 4115 14716
rect 3819 14662 3865 14714
rect 3865 14662 3875 14714
rect 3899 14662 3929 14714
rect 3929 14662 3941 14714
rect 3941 14662 3955 14714
rect 3979 14662 3993 14714
rect 3993 14662 4005 14714
rect 4005 14662 4035 14714
rect 4059 14662 4069 14714
rect 4069 14662 4115 14714
rect 3819 14660 3875 14662
rect 3899 14660 3955 14662
rect 3979 14660 4035 14662
rect 4059 14660 4115 14662
rect 846 14456 902 14512
rect 4479 14170 4535 14172
rect 4559 14170 4615 14172
rect 4639 14170 4695 14172
rect 4719 14170 4775 14172
rect 4479 14118 4525 14170
rect 4525 14118 4535 14170
rect 4559 14118 4589 14170
rect 4589 14118 4601 14170
rect 4601 14118 4615 14170
rect 4639 14118 4653 14170
rect 4653 14118 4665 14170
rect 4665 14118 4695 14170
rect 4719 14118 4729 14170
rect 4729 14118 4775 14170
rect 4479 14116 4535 14118
rect 4559 14116 4615 14118
rect 4639 14116 4695 14118
rect 4719 14116 4775 14118
rect 1398 13640 1454 13696
rect 3819 13626 3875 13628
rect 3899 13626 3955 13628
rect 3979 13626 4035 13628
rect 4059 13626 4115 13628
rect 3819 13574 3865 13626
rect 3865 13574 3875 13626
rect 3899 13574 3929 13626
rect 3929 13574 3941 13626
rect 3941 13574 3955 13626
rect 3979 13574 3993 13626
rect 3993 13574 4005 13626
rect 4005 13574 4035 13626
rect 4059 13574 4069 13626
rect 4069 13574 4115 13626
rect 3819 13572 3875 13574
rect 3899 13572 3955 13574
rect 3979 13572 4035 13574
rect 4059 13572 4115 13574
rect 846 13096 902 13152
rect 4479 13082 4535 13084
rect 4559 13082 4615 13084
rect 4639 13082 4695 13084
rect 4719 13082 4775 13084
rect 4479 13030 4525 13082
rect 4525 13030 4535 13082
rect 4559 13030 4589 13082
rect 4589 13030 4601 13082
rect 4601 13030 4615 13082
rect 4639 13030 4653 13082
rect 4653 13030 4665 13082
rect 4665 13030 4695 13082
rect 4719 13030 4729 13082
rect 4729 13030 4775 13082
rect 4479 13028 4535 13030
rect 4559 13028 4615 13030
rect 4639 13028 4695 13030
rect 4719 13028 4775 13030
rect 3819 12538 3875 12540
rect 3899 12538 3955 12540
rect 3979 12538 4035 12540
rect 4059 12538 4115 12540
rect 3819 12486 3865 12538
rect 3865 12486 3875 12538
rect 3899 12486 3929 12538
rect 3929 12486 3941 12538
rect 3941 12486 3955 12538
rect 3979 12486 3993 12538
rect 3993 12486 4005 12538
rect 4005 12486 4035 12538
rect 4059 12486 4069 12538
rect 4069 12486 4115 12538
rect 3819 12484 3875 12486
rect 3899 12484 3955 12486
rect 3979 12484 4035 12486
rect 4059 12484 4115 12486
rect 1398 12280 1454 12336
rect 846 11756 902 11792
rect 9546 17978 9602 17980
rect 9626 17978 9682 17980
rect 9706 17978 9762 17980
rect 9786 17978 9842 17980
rect 9546 17926 9592 17978
rect 9592 17926 9602 17978
rect 9626 17926 9656 17978
rect 9656 17926 9668 17978
rect 9668 17926 9682 17978
rect 9706 17926 9720 17978
rect 9720 17926 9732 17978
rect 9732 17926 9762 17978
rect 9786 17926 9796 17978
rect 9796 17926 9842 17978
rect 9546 17924 9602 17926
rect 9626 17924 9682 17926
rect 9706 17924 9762 17926
rect 9786 17924 9842 17926
rect 10206 23962 10262 23964
rect 10286 23962 10342 23964
rect 10366 23962 10422 23964
rect 10446 23962 10502 23964
rect 10206 23910 10252 23962
rect 10252 23910 10262 23962
rect 10286 23910 10316 23962
rect 10316 23910 10328 23962
rect 10328 23910 10342 23962
rect 10366 23910 10380 23962
rect 10380 23910 10392 23962
rect 10392 23910 10422 23962
rect 10446 23910 10456 23962
rect 10456 23910 10502 23962
rect 10206 23908 10262 23910
rect 10286 23908 10342 23910
rect 10366 23908 10422 23910
rect 10446 23908 10502 23910
rect 10206 22874 10262 22876
rect 10286 22874 10342 22876
rect 10366 22874 10422 22876
rect 10446 22874 10502 22876
rect 10206 22822 10252 22874
rect 10252 22822 10262 22874
rect 10286 22822 10316 22874
rect 10316 22822 10328 22874
rect 10328 22822 10342 22874
rect 10366 22822 10380 22874
rect 10380 22822 10392 22874
rect 10392 22822 10422 22874
rect 10446 22822 10456 22874
rect 10456 22822 10502 22874
rect 10206 22820 10262 22822
rect 10286 22820 10342 22822
rect 10366 22820 10422 22822
rect 10446 22820 10502 22822
rect 10206 21786 10262 21788
rect 10286 21786 10342 21788
rect 10366 21786 10422 21788
rect 10446 21786 10502 21788
rect 10206 21734 10252 21786
rect 10252 21734 10262 21786
rect 10286 21734 10316 21786
rect 10316 21734 10328 21786
rect 10328 21734 10342 21786
rect 10366 21734 10380 21786
rect 10380 21734 10392 21786
rect 10392 21734 10422 21786
rect 10446 21734 10456 21786
rect 10456 21734 10502 21786
rect 10206 21732 10262 21734
rect 10286 21732 10342 21734
rect 10366 21732 10422 21734
rect 10446 21732 10502 21734
rect 10206 20698 10262 20700
rect 10286 20698 10342 20700
rect 10366 20698 10422 20700
rect 10446 20698 10502 20700
rect 10206 20646 10252 20698
rect 10252 20646 10262 20698
rect 10286 20646 10316 20698
rect 10316 20646 10328 20698
rect 10328 20646 10342 20698
rect 10366 20646 10380 20698
rect 10380 20646 10392 20698
rect 10392 20646 10422 20698
rect 10446 20646 10456 20698
rect 10456 20646 10502 20698
rect 10206 20644 10262 20646
rect 10286 20644 10342 20646
rect 10366 20644 10422 20646
rect 10446 20644 10502 20646
rect 10206 19610 10262 19612
rect 10286 19610 10342 19612
rect 10366 19610 10422 19612
rect 10446 19610 10502 19612
rect 10206 19558 10252 19610
rect 10252 19558 10262 19610
rect 10286 19558 10316 19610
rect 10316 19558 10328 19610
rect 10328 19558 10342 19610
rect 10366 19558 10380 19610
rect 10380 19558 10392 19610
rect 10392 19558 10422 19610
rect 10446 19558 10456 19610
rect 10456 19558 10502 19610
rect 10206 19556 10262 19558
rect 10286 19556 10342 19558
rect 10366 19556 10422 19558
rect 10446 19556 10502 19558
rect 10206 18522 10262 18524
rect 10286 18522 10342 18524
rect 10366 18522 10422 18524
rect 10446 18522 10502 18524
rect 10206 18470 10252 18522
rect 10252 18470 10262 18522
rect 10286 18470 10316 18522
rect 10316 18470 10328 18522
rect 10328 18470 10342 18522
rect 10366 18470 10380 18522
rect 10380 18470 10392 18522
rect 10392 18470 10422 18522
rect 10446 18470 10456 18522
rect 10456 18470 10502 18522
rect 10206 18468 10262 18470
rect 10286 18468 10342 18470
rect 10366 18468 10422 18470
rect 10446 18468 10502 18470
rect 10206 17434 10262 17436
rect 10286 17434 10342 17436
rect 10366 17434 10422 17436
rect 10446 17434 10502 17436
rect 10206 17382 10252 17434
rect 10252 17382 10262 17434
rect 10286 17382 10316 17434
rect 10316 17382 10328 17434
rect 10328 17382 10342 17434
rect 10366 17382 10380 17434
rect 10380 17382 10392 17434
rect 10392 17382 10422 17434
rect 10446 17382 10456 17434
rect 10456 17382 10502 17434
rect 10206 17380 10262 17382
rect 10286 17380 10342 17382
rect 10366 17380 10422 17382
rect 10446 17380 10502 17382
rect 9546 16890 9602 16892
rect 9626 16890 9682 16892
rect 9706 16890 9762 16892
rect 9786 16890 9842 16892
rect 9546 16838 9592 16890
rect 9592 16838 9602 16890
rect 9626 16838 9656 16890
rect 9656 16838 9668 16890
rect 9668 16838 9682 16890
rect 9706 16838 9720 16890
rect 9720 16838 9732 16890
rect 9732 16838 9762 16890
rect 9786 16838 9796 16890
rect 9796 16838 9842 16890
rect 9546 16836 9602 16838
rect 9626 16836 9682 16838
rect 9706 16836 9762 16838
rect 9786 16836 9842 16838
rect 4479 11994 4535 11996
rect 4559 11994 4615 11996
rect 4639 11994 4695 11996
rect 4719 11994 4775 11996
rect 4479 11942 4525 11994
rect 4525 11942 4535 11994
rect 4559 11942 4589 11994
rect 4589 11942 4601 11994
rect 4601 11942 4615 11994
rect 4639 11942 4653 11994
rect 4653 11942 4665 11994
rect 4665 11942 4695 11994
rect 4719 11942 4729 11994
rect 4729 11942 4775 11994
rect 4479 11940 4535 11942
rect 4559 11940 4615 11942
rect 4639 11940 4695 11942
rect 4719 11940 4775 11942
rect 846 11736 848 11756
rect 848 11736 900 11756
rect 900 11736 902 11756
rect 3819 11450 3875 11452
rect 3899 11450 3955 11452
rect 3979 11450 4035 11452
rect 4059 11450 4115 11452
rect 3819 11398 3865 11450
rect 3865 11398 3875 11450
rect 3899 11398 3929 11450
rect 3929 11398 3941 11450
rect 3941 11398 3955 11450
rect 3979 11398 3993 11450
rect 3993 11398 4005 11450
rect 4005 11398 4035 11450
rect 4059 11398 4069 11450
rect 4069 11398 4115 11450
rect 3819 11396 3875 11398
rect 3899 11396 3955 11398
rect 3979 11396 4035 11398
rect 4059 11396 4115 11398
rect 1398 10920 1454 10976
rect 4479 10906 4535 10908
rect 4559 10906 4615 10908
rect 4639 10906 4695 10908
rect 4719 10906 4775 10908
rect 4479 10854 4525 10906
rect 4525 10854 4535 10906
rect 4559 10854 4589 10906
rect 4589 10854 4601 10906
rect 4601 10854 4615 10906
rect 4639 10854 4653 10906
rect 4653 10854 4665 10906
rect 4665 10854 4695 10906
rect 4719 10854 4729 10906
rect 4729 10854 4775 10906
rect 4479 10852 4535 10854
rect 4559 10852 4615 10854
rect 4639 10852 4695 10854
rect 4719 10852 4775 10854
rect 846 10412 848 10432
rect 848 10412 900 10432
rect 900 10412 902 10432
rect 846 10376 902 10412
rect 3819 10362 3875 10364
rect 3899 10362 3955 10364
rect 3979 10362 4035 10364
rect 4059 10362 4115 10364
rect 3819 10310 3865 10362
rect 3865 10310 3875 10362
rect 3899 10310 3929 10362
rect 3929 10310 3941 10362
rect 3941 10310 3955 10362
rect 3979 10310 3993 10362
rect 3993 10310 4005 10362
rect 4005 10310 4035 10362
rect 4059 10310 4069 10362
rect 4069 10310 4115 10362
rect 3819 10308 3875 10310
rect 3899 10308 3955 10310
rect 3979 10308 4035 10310
rect 4059 10308 4115 10310
rect 4479 9818 4535 9820
rect 4559 9818 4615 9820
rect 4639 9818 4695 9820
rect 4719 9818 4775 9820
rect 4479 9766 4525 9818
rect 4525 9766 4535 9818
rect 4559 9766 4589 9818
rect 4589 9766 4601 9818
rect 4601 9766 4615 9818
rect 4639 9766 4653 9818
rect 4653 9766 4665 9818
rect 4665 9766 4695 9818
rect 4719 9766 4729 9818
rect 4729 9766 4775 9818
rect 4479 9764 4535 9766
rect 4559 9764 4615 9766
rect 4639 9764 4695 9766
rect 4719 9764 4775 9766
rect 1398 9560 1454 9616
rect 3819 9274 3875 9276
rect 3899 9274 3955 9276
rect 3979 9274 4035 9276
rect 4059 9274 4115 9276
rect 3819 9222 3865 9274
rect 3865 9222 3875 9274
rect 3899 9222 3929 9274
rect 3929 9222 3941 9274
rect 3941 9222 3955 9274
rect 3979 9222 3993 9274
rect 3993 9222 4005 9274
rect 4005 9222 4035 9274
rect 4059 9222 4069 9274
rect 4069 9222 4115 9274
rect 3819 9220 3875 9222
rect 3899 9220 3955 9222
rect 3979 9220 4035 9222
rect 4059 9220 4115 9222
rect 846 9052 848 9072
rect 848 9052 900 9072
rect 900 9052 902 9072
rect 846 9016 902 9052
rect 4479 8730 4535 8732
rect 4559 8730 4615 8732
rect 4639 8730 4695 8732
rect 4719 8730 4775 8732
rect 4479 8678 4525 8730
rect 4525 8678 4535 8730
rect 4559 8678 4589 8730
rect 4589 8678 4601 8730
rect 4601 8678 4615 8730
rect 4639 8678 4653 8730
rect 4653 8678 4665 8730
rect 4665 8678 4695 8730
rect 4719 8678 4729 8730
rect 4729 8678 4775 8730
rect 4479 8676 4535 8678
rect 4559 8676 4615 8678
rect 4639 8676 4695 8678
rect 4719 8676 4775 8678
rect 3819 8186 3875 8188
rect 3899 8186 3955 8188
rect 3979 8186 4035 8188
rect 4059 8186 4115 8188
rect 3819 8134 3865 8186
rect 3865 8134 3875 8186
rect 3899 8134 3929 8186
rect 3929 8134 3941 8186
rect 3941 8134 3955 8186
rect 3979 8134 3993 8186
rect 3993 8134 4005 8186
rect 4005 8134 4035 8186
rect 4059 8134 4069 8186
rect 4069 8134 4115 8186
rect 3819 8132 3875 8134
rect 3899 8132 3955 8134
rect 3979 8132 4035 8134
rect 4059 8132 4115 8134
rect 846 7656 902 7712
rect 4479 7642 4535 7644
rect 4559 7642 4615 7644
rect 4639 7642 4695 7644
rect 4719 7642 4775 7644
rect 4479 7590 4525 7642
rect 4525 7590 4535 7642
rect 4559 7590 4589 7642
rect 4589 7590 4601 7642
rect 4601 7590 4615 7642
rect 4639 7590 4653 7642
rect 4653 7590 4665 7642
rect 4665 7590 4695 7642
rect 4719 7590 4729 7642
rect 4729 7590 4775 7642
rect 4479 7588 4535 7590
rect 4559 7588 4615 7590
rect 4639 7588 4695 7590
rect 4719 7588 4775 7590
rect 3819 7098 3875 7100
rect 3899 7098 3955 7100
rect 3979 7098 4035 7100
rect 4059 7098 4115 7100
rect 3819 7046 3865 7098
rect 3865 7046 3875 7098
rect 3899 7046 3929 7098
rect 3929 7046 3941 7098
rect 3941 7046 3955 7098
rect 3979 7046 3993 7098
rect 3993 7046 4005 7098
rect 4005 7046 4035 7098
rect 4059 7046 4069 7098
rect 4069 7046 4115 7098
rect 3819 7044 3875 7046
rect 3899 7044 3955 7046
rect 3979 7044 4035 7046
rect 4059 7044 4115 7046
rect 1398 6840 1454 6896
rect 3819 6010 3875 6012
rect 3899 6010 3955 6012
rect 3979 6010 4035 6012
rect 4059 6010 4115 6012
rect 3819 5958 3865 6010
rect 3865 5958 3875 6010
rect 3899 5958 3929 6010
rect 3929 5958 3941 6010
rect 3941 5958 3955 6010
rect 3979 5958 3993 6010
rect 3993 5958 4005 6010
rect 4005 5958 4035 6010
rect 4059 5958 4069 6010
rect 4069 5958 4115 6010
rect 3819 5956 3875 5958
rect 3899 5956 3955 5958
rect 3979 5956 4035 5958
rect 4059 5956 4115 5958
rect 3819 4922 3875 4924
rect 3899 4922 3955 4924
rect 3979 4922 4035 4924
rect 4059 4922 4115 4924
rect 3819 4870 3865 4922
rect 3865 4870 3875 4922
rect 3899 4870 3929 4922
rect 3929 4870 3941 4922
rect 3941 4870 3955 4922
rect 3979 4870 3993 4922
rect 3993 4870 4005 4922
rect 4005 4870 4035 4922
rect 4059 4870 4069 4922
rect 4069 4870 4115 4922
rect 3819 4868 3875 4870
rect 3899 4868 3955 4870
rect 3979 4868 4035 4870
rect 4059 4868 4115 4870
rect 3819 3834 3875 3836
rect 3899 3834 3955 3836
rect 3979 3834 4035 3836
rect 4059 3834 4115 3836
rect 3819 3782 3865 3834
rect 3865 3782 3875 3834
rect 3899 3782 3929 3834
rect 3929 3782 3941 3834
rect 3941 3782 3955 3834
rect 3979 3782 3993 3834
rect 3993 3782 4005 3834
rect 4005 3782 4035 3834
rect 4059 3782 4069 3834
rect 4069 3782 4115 3834
rect 3819 3780 3875 3782
rect 3899 3780 3955 3782
rect 3979 3780 4035 3782
rect 4059 3780 4115 3782
rect 3819 2746 3875 2748
rect 3899 2746 3955 2748
rect 3979 2746 4035 2748
rect 4059 2746 4115 2748
rect 3819 2694 3865 2746
rect 3865 2694 3875 2746
rect 3899 2694 3929 2746
rect 3929 2694 3941 2746
rect 3941 2694 3955 2746
rect 3979 2694 3993 2746
rect 3993 2694 4005 2746
rect 4005 2694 4035 2746
rect 4059 2694 4069 2746
rect 4069 2694 4115 2746
rect 3819 2692 3875 2694
rect 3899 2692 3955 2694
rect 3979 2692 4035 2694
rect 4059 2692 4115 2694
rect 4479 6554 4535 6556
rect 4559 6554 4615 6556
rect 4639 6554 4695 6556
rect 4719 6554 4775 6556
rect 4479 6502 4525 6554
rect 4525 6502 4535 6554
rect 4559 6502 4589 6554
rect 4589 6502 4601 6554
rect 4601 6502 4615 6554
rect 4639 6502 4653 6554
rect 4653 6502 4665 6554
rect 4665 6502 4695 6554
rect 4719 6502 4729 6554
rect 4729 6502 4775 6554
rect 4479 6500 4535 6502
rect 4559 6500 4615 6502
rect 4639 6500 4695 6502
rect 4719 6500 4775 6502
rect 4479 5466 4535 5468
rect 4559 5466 4615 5468
rect 4639 5466 4695 5468
rect 4719 5466 4775 5468
rect 4479 5414 4525 5466
rect 4525 5414 4535 5466
rect 4559 5414 4589 5466
rect 4589 5414 4601 5466
rect 4601 5414 4615 5466
rect 4639 5414 4653 5466
rect 4653 5414 4665 5466
rect 4665 5414 4695 5466
rect 4719 5414 4729 5466
rect 4729 5414 4775 5466
rect 4479 5412 4535 5414
rect 4559 5412 4615 5414
rect 4639 5412 4695 5414
rect 4719 5412 4775 5414
rect 4479 4378 4535 4380
rect 4559 4378 4615 4380
rect 4639 4378 4695 4380
rect 4719 4378 4775 4380
rect 4479 4326 4525 4378
rect 4525 4326 4535 4378
rect 4559 4326 4589 4378
rect 4589 4326 4601 4378
rect 4601 4326 4615 4378
rect 4639 4326 4653 4378
rect 4653 4326 4665 4378
rect 4665 4326 4695 4378
rect 4719 4326 4729 4378
rect 4729 4326 4775 4378
rect 4479 4324 4535 4326
rect 4559 4324 4615 4326
rect 4639 4324 4695 4326
rect 4719 4324 4775 4326
rect 10206 16346 10262 16348
rect 10286 16346 10342 16348
rect 10366 16346 10422 16348
rect 10446 16346 10502 16348
rect 10206 16294 10252 16346
rect 10252 16294 10262 16346
rect 10286 16294 10316 16346
rect 10316 16294 10328 16346
rect 10328 16294 10342 16346
rect 10366 16294 10380 16346
rect 10380 16294 10392 16346
rect 10392 16294 10422 16346
rect 10446 16294 10456 16346
rect 10456 16294 10502 16346
rect 10206 16292 10262 16294
rect 10286 16292 10342 16294
rect 10366 16292 10422 16294
rect 10446 16292 10502 16294
rect 9546 15802 9602 15804
rect 9626 15802 9682 15804
rect 9706 15802 9762 15804
rect 9786 15802 9842 15804
rect 9546 15750 9592 15802
rect 9592 15750 9602 15802
rect 9626 15750 9656 15802
rect 9656 15750 9668 15802
rect 9668 15750 9682 15802
rect 9706 15750 9720 15802
rect 9720 15750 9732 15802
rect 9732 15750 9762 15802
rect 9786 15750 9796 15802
rect 9796 15750 9842 15802
rect 9546 15748 9602 15750
rect 9626 15748 9682 15750
rect 9706 15748 9762 15750
rect 9786 15748 9842 15750
rect 9546 14714 9602 14716
rect 9626 14714 9682 14716
rect 9706 14714 9762 14716
rect 9786 14714 9842 14716
rect 9546 14662 9592 14714
rect 9592 14662 9602 14714
rect 9626 14662 9656 14714
rect 9656 14662 9668 14714
rect 9668 14662 9682 14714
rect 9706 14662 9720 14714
rect 9720 14662 9732 14714
rect 9732 14662 9762 14714
rect 9786 14662 9796 14714
rect 9796 14662 9842 14714
rect 9546 14660 9602 14662
rect 9626 14660 9682 14662
rect 9706 14660 9762 14662
rect 9786 14660 9842 14662
rect 10206 15258 10262 15260
rect 10286 15258 10342 15260
rect 10366 15258 10422 15260
rect 10446 15258 10502 15260
rect 10206 15206 10252 15258
rect 10252 15206 10262 15258
rect 10286 15206 10316 15258
rect 10316 15206 10328 15258
rect 10328 15206 10342 15258
rect 10366 15206 10380 15258
rect 10380 15206 10392 15258
rect 10392 15206 10422 15258
rect 10446 15206 10456 15258
rect 10456 15206 10502 15258
rect 10206 15204 10262 15206
rect 10286 15204 10342 15206
rect 10366 15204 10422 15206
rect 10446 15204 10502 15206
rect 9546 13626 9602 13628
rect 9626 13626 9682 13628
rect 9706 13626 9762 13628
rect 9786 13626 9842 13628
rect 9546 13574 9592 13626
rect 9592 13574 9602 13626
rect 9626 13574 9656 13626
rect 9656 13574 9668 13626
rect 9668 13574 9682 13626
rect 9706 13574 9720 13626
rect 9720 13574 9732 13626
rect 9732 13574 9762 13626
rect 9786 13574 9796 13626
rect 9796 13574 9842 13626
rect 9546 13572 9602 13574
rect 9626 13572 9682 13574
rect 9706 13572 9762 13574
rect 9786 13572 9842 13574
rect 10206 14170 10262 14172
rect 10286 14170 10342 14172
rect 10366 14170 10422 14172
rect 10446 14170 10502 14172
rect 10206 14118 10252 14170
rect 10252 14118 10262 14170
rect 10286 14118 10316 14170
rect 10316 14118 10328 14170
rect 10328 14118 10342 14170
rect 10366 14118 10380 14170
rect 10380 14118 10392 14170
rect 10392 14118 10422 14170
rect 10446 14118 10456 14170
rect 10456 14118 10502 14170
rect 10206 14116 10262 14118
rect 10286 14116 10342 14118
rect 10366 14116 10422 14118
rect 10446 14116 10502 14118
rect 10206 13082 10262 13084
rect 10286 13082 10342 13084
rect 10366 13082 10422 13084
rect 10446 13082 10502 13084
rect 10206 13030 10252 13082
rect 10252 13030 10262 13082
rect 10286 13030 10316 13082
rect 10316 13030 10328 13082
rect 10328 13030 10342 13082
rect 10366 13030 10380 13082
rect 10380 13030 10392 13082
rect 10392 13030 10422 13082
rect 10446 13030 10456 13082
rect 10456 13030 10502 13082
rect 10206 13028 10262 13030
rect 10286 13028 10342 13030
rect 10366 13028 10422 13030
rect 10446 13028 10502 13030
rect 9546 12538 9602 12540
rect 9626 12538 9682 12540
rect 9706 12538 9762 12540
rect 9786 12538 9842 12540
rect 9546 12486 9592 12538
rect 9592 12486 9602 12538
rect 9626 12486 9656 12538
rect 9656 12486 9668 12538
rect 9668 12486 9682 12538
rect 9706 12486 9720 12538
rect 9720 12486 9732 12538
rect 9732 12486 9762 12538
rect 9786 12486 9796 12538
rect 9796 12486 9842 12538
rect 9546 12484 9602 12486
rect 9626 12484 9682 12486
rect 9706 12484 9762 12486
rect 9786 12484 9842 12486
rect 10206 11994 10262 11996
rect 10286 11994 10342 11996
rect 10366 11994 10422 11996
rect 10446 11994 10502 11996
rect 10206 11942 10252 11994
rect 10252 11942 10262 11994
rect 10286 11942 10316 11994
rect 10316 11942 10328 11994
rect 10328 11942 10342 11994
rect 10366 11942 10380 11994
rect 10380 11942 10392 11994
rect 10392 11942 10422 11994
rect 10446 11942 10456 11994
rect 10456 11942 10502 11994
rect 10206 11940 10262 11942
rect 10286 11940 10342 11942
rect 10366 11940 10422 11942
rect 10446 11940 10502 11942
rect 9546 11450 9602 11452
rect 9626 11450 9682 11452
rect 9706 11450 9762 11452
rect 9786 11450 9842 11452
rect 9546 11398 9592 11450
rect 9592 11398 9602 11450
rect 9626 11398 9656 11450
rect 9656 11398 9668 11450
rect 9668 11398 9682 11450
rect 9706 11398 9720 11450
rect 9720 11398 9732 11450
rect 9732 11398 9762 11450
rect 9786 11398 9796 11450
rect 9796 11398 9842 11450
rect 9546 11396 9602 11398
rect 9626 11396 9682 11398
rect 9706 11396 9762 11398
rect 9786 11396 9842 11398
rect 4479 3290 4535 3292
rect 4559 3290 4615 3292
rect 4639 3290 4695 3292
rect 4719 3290 4775 3292
rect 4479 3238 4525 3290
rect 4525 3238 4535 3290
rect 4559 3238 4589 3290
rect 4589 3238 4601 3290
rect 4601 3238 4615 3290
rect 4639 3238 4653 3290
rect 4653 3238 4665 3290
rect 4665 3238 4695 3290
rect 4719 3238 4729 3290
rect 4729 3238 4775 3290
rect 4479 3236 4535 3238
rect 4559 3236 4615 3238
rect 4639 3236 4695 3238
rect 4719 3236 4775 3238
rect 10206 10906 10262 10908
rect 10286 10906 10342 10908
rect 10366 10906 10422 10908
rect 10446 10906 10502 10908
rect 10206 10854 10252 10906
rect 10252 10854 10262 10906
rect 10286 10854 10316 10906
rect 10316 10854 10328 10906
rect 10328 10854 10342 10906
rect 10366 10854 10380 10906
rect 10380 10854 10392 10906
rect 10392 10854 10422 10906
rect 10446 10854 10456 10906
rect 10456 10854 10502 10906
rect 10206 10852 10262 10854
rect 10286 10852 10342 10854
rect 10366 10852 10422 10854
rect 10446 10852 10502 10854
rect 9546 10362 9602 10364
rect 9626 10362 9682 10364
rect 9706 10362 9762 10364
rect 9786 10362 9842 10364
rect 9546 10310 9592 10362
rect 9592 10310 9602 10362
rect 9626 10310 9656 10362
rect 9656 10310 9668 10362
rect 9668 10310 9682 10362
rect 9706 10310 9720 10362
rect 9720 10310 9732 10362
rect 9732 10310 9762 10362
rect 9786 10310 9796 10362
rect 9796 10310 9842 10362
rect 9546 10308 9602 10310
rect 9626 10308 9682 10310
rect 9706 10308 9762 10310
rect 9786 10308 9842 10310
rect 10206 9818 10262 9820
rect 10286 9818 10342 9820
rect 10366 9818 10422 9820
rect 10446 9818 10502 9820
rect 10206 9766 10252 9818
rect 10252 9766 10262 9818
rect 10286 9766 10316 9818
rect 10316 9766 10328 9818
rect 10328 9766 10342 9818
rect 10366 9766 10380 9818
rect 10380 9766 10392 9818
rect 10392 9766 10422 9818
rect 10446 9766 10456 9818
rect 10456 9766 10502 9818
rect 10206 9764 10262 9766
rect 10286 9764 10342 9766
rect 10366 9764 10422 9766
rect 10446 9764 10502 9766
rect 9546 9274 9602 9276
rect 9626 9274 9682 9276
rect 9706 9274 9762 9276
rect 9786 9274 9842 9276
rect 9546 9222 9592 9274
rect 9592 9222 9602 9274
rect 9626 9222 9656 9274
rect 9656 9222 9668 9274
rect 9668 9222 9682 9274
rect 9706 9222 9720 9274
rect 9720 9222 9732 9274
rect 9732 9222 9762 9274
rect 9786 9222 9796 9274
rect 9796 9222 9842 9274
rect 9546 9220 9602 9222
rect 9626 9220 9682 9222
rect 9706 9220 9762 9222
rect 9786 9220 9842 9222
rect 10206 8730 10262 8732
rect 10286 8730 10342 8732
rect 10366 8730 10422 8732
rect 10446 8730 10502 8732
rect 10206 8678 10252 8730
rect 10252 8678 10262 8730
rect 10286 8678 10316 8730
rect 10316 8678 10328 8730
rect 10328 8678 10342 8730
rect 10366 8678 10380 8730
rect 10380 8678 10392 8730
rect 10392 8678 10422 8730
rect 10446 8678 10456 8730
rect 10456 8678 10502 8730
rect 10206 8676 10262 8678
rect 10286 8676 10342 8678
rect 10366 8676 10422 8678
rect 10446 8676 10502 8678
rect 9546 8186 9602 8188
rect 9626 8186 9682 8188
rect 9706 8186 9762 8188
rect 9786 8186 9842 8188
rect 9546 8134 9592 8186
rect 9592 8134 9602 8186
rect 9626 8134 9656 8186
rect 9656 8134 9668 8186
rect 9668 8134 9682 8186
rect 9706 8134 9720 8186
rect 9720 8134 9732 8186
rect 9732 8134 9762 8186
rect 9786 8134 9796 8186
rect 9796 8134 9842 8186
rect 9546 8132 9602 8134
rect 9626 8132 9682 8134
rect 9706 8132 9762 8134
rect 9786 8132 9842 8134
rect 10206 7642 10262 7644
rect 10286 7642 10342 7644
rect 10366 7642 10422 7644
rect 10446 7642 10502 7644
rect 10206 7590 10252 7642
rect 10252 7590 10262 7642
rect 10286 7590 10316 7642
rect 10316 7590 10328 7642
rect 10328 7590 10342 7642
rect 10366 7590 10380 7642
rect 10380 7590 10392 7642
rect 10392 7590 10422 7642
rect 10446 7590 10456 7642
rect 10456 7590 10502 7642
rect 10206 7588 10262 7590
rect 10286 7588 10342 7590
rect 10366 7588 10422 7590
rect 10446 7588 10502 7590
rect 9546 7098 9602 7100
rect 9626 7098 9682 7100
rect 9706 7098 9762 7100
rect 9786 7098 9842 7100
rect 9546 7046 9592 7098
rect 9592 7046 9602 7098
rect 9626 7046 9656 7098
rect 9656 7046 9668 7098
rect 9668 7046 9682 7098
rect 9706 7046 9720 7098
rect 9720 7046 9732 7098
rect 9732 7046 9762 7098
rect 9786 7046 9796 7098
rect 9796 7046 9842 7098
rect 9546 7044 9602 7046
rect 9626 7044 9682 7046
rect 9706 7044 9762 7046
rect 9786 7044 9842 7046
rect 9546 6010 9602 6012
rect 9626 6010 9682 6012
rect 9706 6010 9762 6012
rect 9786 6010 9842 6012
rect 9546 5958 9592 6010
rect 9592 5958 9602 6010
rect 9626 5958 9656 6010
rect 9656 5958 9668 6010
rect 9668 5958 9682 6010
rect 9706 5958 9720 6010
rect 9720 5958 9732 6010
rect 9732 5958 9762 6010
rect 9786 5958 9796 6010
rect 9796 5958 9842 6010
rect 9546 5956 9602 5958
rect 9626 5956 9682 5958
rect 9706 5956 9762 5958
rect 9786 5956 9842 5958
rect 9546 4922 9602 4924
rect 9626 4922 9682 4924
rect 9706 4922 9762 4924
rect 9786 4922 9842 4924
rect 9546 4870 9592 4922
rect 9592 4870 9602 4922
rect 9626 4870 9656 4922
rect 9656 4870 9668 4922
rect 9668 4870 9682 4922
rect 9706 4870 9720 4922
rect 9720 4870 9732 4922
rect 9732 4870 9762 4922
rect 9786 4870 9796 4922
rect 9796 4870 9842 4922
rect 9546 4868 9602 4870
rect 9626 4868 9682 4870
rect 9706 4868 9762 4870
rect 9786 4868 9842 4870
rect 9546 3834 9602 3836
rect 9626 3834 9682 3836
rect 9706 3834 9762 3836
rect 9786 3834 9842 3836
rect 9546 3782 9592 3834
rect 9592 3782 9602 3834
rect 9626 3782 9656 3834
rect 9656 3782 9668 3834
rect 9668 3782 9682 3834
rect 9706 3782 9720 3834
rect 9720 3782 9732 3834
rect 9732 3782 9762 3834
rect 9786 3782 9796 3834
rect 9796 3782 9842 3834
rect 9546 3780 9602 3782
rect 9626 3780 9682 3782
rect 9706 3780 9762 3782
rect 9786 3780 9842 3782
rect 9546 2746 9602 2748
rect 9626 2746 9682 2748
rect 9706 2746 9762 2748
rect 9786 2746 9842 2748
rect 9546 2694 9592 2746
rect 9592 2694 9602 2746
rect 9626 2694 9656 2746
rect 9656 2694 9668 2746
rect 9668 2694 9682 2746
rect 9706 2694 9720 2746
rect 9720 2694 9732 2746
rect 9732 2694 9762 2746
rect 9786 2694 9796 2746
rect 9796 2694 9842 2746
rect 9546 2692 9602 2694
rect 9626 2692 9682 2694
rect 9706 2692 9762 2694
rect 9786 2692 9842 2694
rect 10206 6554 10262 6556
rect 10286 6554 10342 6556
rect 10366 6554 10422 6556
rect 10446 6554 10502 6556
rect 10206 6502 10252 6554
rect 10252 6502 10262 6554
rect 10286 6502 10316 6554
rect 10316 6502 10328 6554
rect 10328 6502 10342 6554
rect 10366 6502 10380 6554
rect 10380 6502 10392 6554
rect 10392 6502 10422 6554
rect 10446 6502 10456 6554
rect 10456 6502 10502 6554
rect 10206 6500 10262 6502
rect 10286 6500 10342 6502
rect 10366 6500 10422 6502
rect 10446 6500 10502 6502
rect 10206 5466 10262 5468
rect 10286 5466 10342 5468
rect 10366 5466 10422 5468
rect 10446 5466 10502 5468
rect 10206 5414 10252 5466
rect 10252 5414 10262 5466
rect 10286 5414 10316 5466
rect 10316 5414 10328 5466
rect 10328 5414 10342 5466
rect 10366 5414 10380 5466
rect 10380 5414 10392 5466
rect 10392 5414 10422 5466
rect 10446 5414 10456 5466
rect 10456 5414 10502 5466
rect 10206 5412 10262 5414
rect 10286 5412 10342 5414
rect 10366 5412 10422 5414
rect 10446 5412 10502 5414
rect 10206 4378 10262 4380
rect 10286 4378 10342 4380
rect 10366 4378 10422 4380
rect 10446 4378 10502 4380
rect 10206 4326 10252 4378
rect 10252 4326 10262 4378
rect 10286 4326 10316 4378
rect 10316 4326 10328 4378
rect 10328 4326 10342 4378
rect 10366 4326 10380 4378
rect 10380 4326 10392 4378
rect 10392 4326 10422 4378
rect 10446 4326 10456 4378
rect 10456 4326 10502 4378
rect 10206 4324 10262 4326
rect 10286 4324 10342 4326
rect 10366 4324 10422 4326
rect 10446 4324 10502 4326
rect 10206 3290 10262 3292
rect 10286 3290 10342 3292
rect 10366 3290 10422 3292
rect 10446 3290 10502 3292
rect 10206 3238 10252 3290
rect 10252 3238 10262 3290
rect 10286 3238 10316 3290
rect 10316 3238 10328 3290
rect 10328 3238 10342 3290
rect 10366 3238 10380 3290
rect 10380 3238 10392 3290
rect 10392 3238 10422 3290
rect 10446 3238 10456 3290
rect 10456 3238 10502 3290
rect 10206 3236 10262 3238
rect 10286 3236 10342 3238
rect 10366 3236 10422 3238
rect 10446 3236 10502 3238
rect 4479 2202 4535 2204
rect 4559 2202 4615 2204
rect 4639 2202 4695 2204
rect 4719 2202 4775 2204
rect 4479 2150 4525 2202
rect 4525 2150 4535 2202
rect 4559 2150 4589 2202
rect 4589 2150 4601 2202
rect 4601 2150 4615 2202
rect 4639 2150 4653 2202
rect 4653 2150 4665 2202
rect 4665 2150 4695 2202
rect 4719 2150 4729 2202
rect 4729 2150 4775 2202
rect 4479 2148 4535 2150
rect 4559 2148 4615 2150
rect 4639 2148 4695 2150
rect 4719 2148 4775 2150
rect 10206 2202 10262 2204
rect 10286 2202 10342 2204
rect 10366 2202 10422 2204
rect 10446 2202 10502 2204
rect 10206 2150 10252 2202
rect 10252 2150 10262 2202
rect 10286 2150 10316 2202
rect 10316 2150 10328 2202
rect 10328 2150 10342 2202
rect 10366 2150 10380 2202
rect 10380 2150 10392 2202
rect 10392 2150 10422 2202
rect 10446 2150 10456 2202
rect 10456 2150 10502 2202
rect 10206 2148 10262 2150
rect 10286 2148 10342 2150
rect 10366 2148 10422 2150
rect 10446 2148 10502 2150
rect 15933 25050 15989 25052
rect 16013 25050 16069 25052
rect 16093 25050 16149 25052
rect 16173 25050 16229 25052
rect 15933 24998 15979 25050
rect 15979 24998 15989 25050
rect 16013 24998 16043 25050
rect 16043 24998 16055 25050
rect 16055 24998 16069 25050
rect 16093 24998 16107 25050
rect 16107 24998 16119 25050
rect 16119 24998 16149 25050
rect 16173 24998 16183 25050
rect 16183 24998 16229 25050
rect 15933 24996 15989 24998
rect 16013 24996 16069 24998
rect 16093 24996 16149 24998
rect 16173 24996 16229 24998
rect 15273 24506 15329 24508
rect 15353 24506 15409 24508
rect 15433 24506 15489 24508
rect 15513 24506 15569 24508
rect 15273 24454 15319 24506
rect 15319 24454 15329 24506
rect 15353 24454 15383 24506
rect 15383 24454 15395 24506
rect 15395 24454 15409 24506
rect 15433 24454 15447 24506
rect 15447 24454 15459 24506
rect 15459 24454 15489 24506
rect 15513 24454 15523 24506
rect 15523 24454 15569 24506
rect 15273 24452 15329 24454
rect 15353 24452 15409 24454
rect 15433 24452 15489 24454
rect 15513 24452 15569 24454
rect 15273 23418 15329 23420
rect 15353 23418 15409 23420
rect 15433 23418 15489 23420
rect 15513 23418 15569 23420
rect 15273 23366 15319 23418
rect 15319 23366 15329 23418
rect 15353 23366 15383 23418
rect 15383 23366 15395 23418
rect 15395 23366 15409 23418
rect 15433 23366 15447 23418
rect 15447 23366 15459 23418
rect 15459 23366 15489 23418
rect 15513 23366 15523 23418
rect 15523 23366 15569 23418
rect 15273 23364 15329 23366
rect 15353 23364 15409 23366
rect 15433 23364 15489 23366
rect 15513 23364 15569 23366
rect 15273 22330 15329 22332
rect 15353 22330 15409 22332
rect 15433 22330 15489 22332
rect 15513 22330 15569 22332
rect 15273 22278 15319 22330
rect 15319 22278 15329 22330
rect 15353 22278 15383 22330
rect 15383 22278 15395 22330
rect 15395 22278 15409 22330
rect 15433 22278 15447 22330
rect 15447 22278 15459 22330
rect 15459 22278 15489 22330
rect 15513 22278 15523 22330
rect 15523 22278 15569 22330
rect 15273 22276 15329 22278
rect 15353 22276 15409 22278
rect 15433 22276 15489 22278
rect 15513 22276 15569 22278
rect 15273 21242 15329 21244
rect 15353 21242 15409 21244
rect 15433 21242 15489 21244
rect 15513 21242 15569 21244
rect 15273 21190 15319 21242
rect 15319 21190 15329 21242
rect 15353 21190 15383 21242
rect 15383 21190 15395 21242
rect 15395 21190 15409 21242
rect 15433 21190 15447 21242
rect 15447 21190 15459 21242
rect 15459 21190 15489 21242
rect 15513 21190 15523 21242
rect 15523 21190 15569 21242
rect 15273 21188 15329 21190
rect 15353 21188 15409 21190
rect 15433 21188 15489 21190
rect 15513 21188 15569 21190
rect 15273 20154 15329 20156
rect 15353 20154 15409 20156
rect 15433 20154 15489 20156
rect 15513 20154 15569 20156
rect 15273 20102 15319 20154
rect 15319 20102 15329 20154
rect 15353 20102 15383 20154
rect 15383 20102 15395 20154
rect 15395 20102 15409 20154
rect 15433 20102 15447 20154
rect 15447 20102 15459 20154
rect 15459 20102 15489 20154
rect 15513 20102 15523 20154
rect 15523 20102 15569 20154
rect 15273 20100 15329 20102
rect 15353 20100 15409 20102
rect 15433 20100 15489 20102
rect 15513 20100 15569 20102
rect 15273 19066 15329 19068
rect 15353 19066 15409 19068
rect 15433 19066 15489 19068
rect 15513 19066 15569 19068
rect 15273 19014 15319 19066
rect 15319 19014 15329 19066
rect 15353 19014 15383 19066
rect 15383 19014 15395 19066
rect 15395 19014 15409 19066
rect 15433 19014 15447 19066
rect 15447 19014 15459 19066
rect 15459 19014 15489 19066
rect 15513 19014 15523 19066
rect 15523 19014 15569 19066
rect 15273 19012 15329 19014
rect 15353 19012 15409 19014
rect 15433 19012 15489 19014
rect 15513 19012 15569 19014
rect 15273 17978 15329 17980
rect 15353 17978 15409 17980
rect 15433 17978 15489 17980
rect 15513 17978 15569 17980
rect 15273 17926 15319 17978
rect 15319 17926 15329 17978
rect 15353 17926 15383 17978
rect 15383 17926 15395 17978
rect 15395 17926 15409 17978
rect 15433 17926 15447 17978
rect 15447 17926 15459 17978
rect 15459 17926 15489 17978
rect 15513 17926 15523 17978
rect 15523 17926 15569 17978
rect 15273 17924 15329 17926
rect 15353 17924 15409 17926
rect 15433 17924 15489 17926
rect 15513 17924 15569 17926
rect 15273 16890 15329 16892
rect 15353 16890 15409 16892
rect 15433 16890 15489 16892
rect 15513 16890 15569 16892
rect 15273 16838 15319 16890
rect 15319 16838 15329 16890
rect 15353 16838 15383 16890
rect 15383 16838 15395 16890
rect 15395 16838 15409 16890
rect 15433 16838 15447 16890
rect 15447 16838 15459 16890
rect 15459 16838 15489 16890
rect 15513 16838 15523 16890
rect 15523 16838 15569 16890
rect 15273 16836 15329 16838
rect 15353 16836 15409 16838
rect 15433 16836 15489 16838
rect 15513 16836 15569 16838
rect 21660 25050 21716 25052
rect 21740 25050 21796 25052
rect 21820 25050 21876 25052
rect 21900 25050 21956 25052
rect 21660 24998 21706 25050
rect 21706 24998 21716 25050
rect 21740 24998 21770 25050
rect 21770 24998 21782 25050
rect 21782 24998 21796 25050
rect 21820 24998 21834 25050
rect 21834 24998 21846 25050
rect 21846 24998 21876 25050
rect 21900 24998 21910 25050
rect 21910 24998 21956 25050
rect 21660 24996 21716 24998
rect 21740 24996 21796 24998
rect 21820 24996 21876 24998
rect 21900 24996 21956 24998
rect 15933 23962 15989 23964
rect 16013 23962 16069 23964
rect 16093 23962 16149 23964
rect 16173 23962 16229 23964
rect 15933 23910 15979 23962
rect 15979 23910 15989 23962
rect 16013 23910 16043 23962
rect 16043 23910 16055 23962
rect 16055 23910 16069 23962
rect 16093 23910 16107 23962
rect 16107 23910 16119 23962
rect 16119 23910 16149 23962
rect 16173 23910 16183 23962
rect 16183 23910 16229 23962
rect 15933 23908 15989 23910
rect 16013 23908 16069 23910
rect 16093 23908 16149 23910
rect 16173 23908 16229 23910
rect 15933 22874 15989 22876
rect 16013 22874 16069 22876
rect 16093 22874 16149 22876
rect 16173 22874 16229 22876
rect 15933 22822 15979 22874
rect 15979 22822 15989 22874
rect 16013 22822 16043 22874
rect 16043 22822 16055 22874
rect 16055 22822 16069 22874
rect 16093 22822 16107 22874
rect 16107 22822 16119 22874
rect 16119 22822 16149 22874
rect 16173 22822 16183 22874
rect 16183 22822 16229 22874
rect 15933 22820 15989 22822
rect 16013 22820 16069 22822
rect 16093 22820 16149 22822
rect 16173 22820 16229 22822
rect 15933 21786 15989 21788
rect 16013 21786 16069 21788
rect 16093 21786 16149 21788
rect 16173 21786 16229 21788
rect 15933 21734 15979 21786
rect 15979 21734 15989 21786
rect 16013 21734 16043 21786
rect 16043 21734 16055 21786
rect 16055 21734 16069 21786
rect 16093 21734 16107 21786
rect 16107 21734 16119 21786
rect 16119 21734 16149 21786
rect 16173 21734 16183 21786
rect 16183 21734 16229 21786
rect 15933 21732 15989 21734
rect 16013 21732 16069 21734
rect 16093 21732 16149 21734
rect 16173 21732 16229 21734
rect 15933 20698 15989 20700
rect 16013 20698 16069 20700
rect 16093 20698 16149 20700
rect 16173 20698 16229 20700
rect 15933 20646 15979 20698
rect 15979 20646 15989 20698
rect 16013 20646 16043 20698
rect 16043 20646 16055 20698
rect 16055 20646 16069 20698
rect 16093 20646 16107 20698
rect 16107 20646 16119 20698
rect 16119 20646 16149 20698
rect 16173 20646 16183 20698
rect 16183 20646 16229 20698
rect 15933 20644 15989 20646
rect 16013 20644 16069 20646
rect 16093 20644 16149 20646
rect 16173 20644 16229 20646
rect 21000 24506 21056 24508
rect 21080 24506 21136 24508
rect 21160 24506 21216 24508
rect 21240 24506 21296 24508
rect 21000 24454 21046 24506
rect 21046 24454 21056 24506
rect 21080 24454 21110 24506
rect 21110 24454 21122 24506
rect 21122 24454 21136 24506
rect 21160 24454 21174 24506
rect 21174 24454 21186 24506
rect 21186 24454 21216 24506
rect 21240 24454 21250 24506
rect 21250 24454 21296 24506
rect 21000 24452 21056 24454
rect 21080 24452 21136 24454
rect 21160 24452 21216 24454
rect 21240 24452 21296 24454
rect 21660 23962 21716 23964
rect 21740 23962 21796 23964
rect 21820 23962 21876 23964
rect 21900 23962 21956 23964
rect 21660 23910 21706 23962
rect 21706 23910 21716 23962
rect 21740 23910 21770 23962
rect 21770 23910 21782 23962
rect 21782 23910 21796 23962
rect 21820 23910 21834 23962
rect 21834 23910 21846 23962
rect 21846 23910 21876 23962
rect 21900 23910 21910 23962
rect 21910 23910 21956 23962
rect 21660 23908 21716 23910
rect 21740 23908 21796 23910
rect 21820 23908 21876 23910
rect 21900 23908 21956 23910
rect 21000 23418 21056 23420
rect 21080 23418 21136 23420
rect 21160 23418 21216 23420
rect 21240 23418 21296 23420
rect 21000 23366 21046 23418
rect 21046 23366 21056 23418
rect 21080 23366 21110 23418
rect 21110 23366 21122 23418
rect 21122 23366 21136 23418
rect 21160 23366 21174 23418
rect 21174 23366 21186 23418
rect 21186 23366 21216 23418
rect 21240 23366 21250 23418
rect 21250 23366 21296 23418
rect 21000 23364 21056 23366
rect 21080 23364 21136 23366
rect 21160 23364 21216 23366
rect 21240 23364 21296 23366
rect 23662 24520 23718 24576
rect 21660 22874 21716 22876
rect 21740 22874 21796 22876
rect 21820 22874 21876 22876
rect 21900 22874 21956 22876
rect 21660 22822 21706 22874
rect 21706 22822 21716 22874
rect 21740 22822 21770 22874
rect 21770 22822 21782 22874
rect 21782 22822 21796 22874
rect 21820 22822 21834 22874
rect 21834 22822 21846 22874
rect 21846 22822 21876 22874
rect 21900 22822 21910 22874
rect 21910 22822 21956 22874
rect 21660 22820 21716 22822
rect 21740 22820 21796 22822
rect 21820 22820 21876 22822
rect 21900 22820 21956 22822
rect 21000 22330 21056 22332
rect 21080 22330 21136 22332
rect 21160 22330 21216 22332
rect 21240 22330 21296 22332
rect 21000 22278 21046 22330
rect 21046 22278 21056 22330
rect 21080 22278 21110 22330
rect 21110 22278 21122 22330
rect 21122 22278 21136 22330
rect 21160 22278 21174 22330
rect 21174 22278 21186 22330
rect 21186 22278 21216 22330
rect 21240 22278 21250 22330
rect 21250 22278 21296 22330
rect 21000 22276 21056 22278
rect 21080 22276 21136 22278
rect 21160 22276 21216 22278
rect 21240 22276 21296 22278
rect 21660 21786 21716 21788
rect 21740 21786 21796 21788
rect 21820 21786 21876 21788
rect 21900 21786 21956 21788
rect 21660 21734 21706 21786
rect 21706 21734 21716 21786
rect 21740 21734 21770 21786
rect 21770 21734 21782 21786
rect 21782 21734 21796 21786
rect 21820 21734 21834 21786
rect 21834 21734 21846 21786
rect 21846 21734 21876 21786
rect 21900 21734 21910 21786
rect 21910 21734 21956 21786
rect 21660 21732 21716 21734
rect 21740 21732 21796 21734
rect 21820 21732 21876 21734
rect 21900 21732 21956 21734
rect 21000 21242 21056 21244
rect 21080 21242 21136 21244
rect 21160 21242 21216 21244
rect 21240 21242 21296 21244
rect 21000 21190 21046 21242
rect 21046 21190 21056 21242
rect 21080 21190 21110 21242
rect 21110 21190 21122 21242
rect 21122 21190 21136 21242
rect 21160 21190 21174 21242
rect 21174 21190 21186 21242
rect 21186 21190 21216 21242
rect 21240 21190 21250 21242
rect 21250 21190 21296 21242
rect 21000 21188 21056 21190
rect 21080 21188 21136 21190
rect 21160 21188 21216 21190
rect 21240 21188 21296 21190
rect 23662 23840 23718 23896
rect 23386 23160 23442 23216
rect 21660 20698 21716 20700
rect 21740 20698 21796 20700
rect 21820 20698 21876 20700
rect 21900 20698 21956 20700
rect 21660 20646 21706 20698
rect 21706 20646 21716 20698
rect 21740 20646 21770 20698
rect 21770 20646 21782 20698
rect 21782 20646 21796 20698
rect 21820 20646 21834 20698
rect 21834 20646 21846 20698
rect 21846 20646 21876 20698
rect 21900 20646 21910 20698
rect 21910 20646 21956 20698
rect 21660 20644 21716 20646
rect 21740 20644 21796 20646
rect 21820 20644 21876 20646
rect 21900 20644 21956 20646
rect 15933 19610 15989 19612
rect 16013 19610 16069 19612
rect 16093 19610 16149 19612
rect 16173 19610 16229 19612
rect 15933 19558 15979 19610
rect 15979 19558 15989 19610
rect 16013 19558 16043 19610
rect 16043 19558 16055 19610
rect 16055 19558 16069 19610
rect 16093 19558 16107 19610
rect 16107 19558 16119 19610
rect 16119 19558 16149 19610
rect 16173 19558 16183 19610
rect 16183 19558 16229 19610
rect 15933 19556 15989 19558
rect 16013 19556 16069 19558
rect 16093 19556 16149 19558
rect 16173 19556 16229 19558
rect 15933 18522 15989 18524
rect 16013 18522 16069 18524
rect 16093 18522 16149 18524
rect 16173 18522 16229 18524
rect 15933 18470 15979 18522
rect 15979 18470 15989 18522
rect 16013 18470 16043 18522
rect 16043 18470 16055 18522
rect 16055 18470 16069 18522
rect 16093 18470 16107 18522
rect 16107 18470 16119 18522
rect 16119 18470 16149 18522
rect 16173 18470 16183 18522
rect 16183 18470 16229 18522
rect 15933 18468 15989 18470
rect 16013 18468 16069 18470
rect 16093 18468 16149 18470
rect 16173 18468 16229 18470
rect 15933 17434 15989 17436
rect 16013 17434 16069 17436
rect 16093 17434 16149 17436
rect 16173 17434 16229 17436
rect 15933 17382 15979 17434
rect 15979 17382 15989 17434
rect 16013 17382 16043 17434
rect 16043 17382 16055 17434
rect 16055 17382 16069 17434
rect 16093 17382 16107 17434
rect 16107 17382 16119 17434
rect 16119 17382 16149 17434
rect 16173 17382 16183 17434
rect 16183 17382 16229 17434
rect 15933 17380 15989 17382
rect 16013 17380 16069 17382
rect 16093 17380 16149 17382
rect 16173 17380 16229 17382
rect 15933 16346 15989 16348
rect 16013 16346 16069 16348
rect 16093 16346 16149 16348
rect 16173 16346 16229 16348
rect 15933 16294 15979 16346
rect 15979 16294 15989 16346
rect 16013 16294 16043 16346
rect 16043 16294 16055 16346
rect 16055 16294 16069 16346
rect 16093 16294 16107 16346
rect 16107 16294 16119 16346
rect 16119 16294 16149 16346
rect 16173 16294 16183 16346
rect 16183 16294 16229 16346
rect 15933 16292 15989 16294
rect 16013 16292 16069 16294
rect 16093 16292 16149 16294
rect 16173 16292 16229 16294
rect 15273 15802 15329 15804
rect 15353 15802 15409 15804
rect 15433 15802 15489 15804
rect 15513 15802 15569 15804
rect 15273 15750 15319 15802
rect 15319 15750 15329 15802
rect 15353 15750 15383 15802
rect 15383 15750 15395 15802
rect 15395 15750 15409 15802
rect 15433 15750 15447 15802
rect 15447 15750 15459 15802
rect 15459 15750 15489 15802
rect 15513 15750 15523 15802
rect 15523 15750 15569 15802
rect 15273 15748 15329 15750
rect 15353 15748 15409 15750
rect 15433 15748 15489 15750
rect 15513 15748 15569 15750
rect 15933 15258 15989 15260
rect 16013 15258 16069 15260
rect 16093 15258 16149 15260
rect 16173 15258 16229 15260
rect 15933 15206 15979 15258
rect 15979 15206 15989 15258
rect 16013 15206 16043 15258
rect 16043 15206 16055 15258
rect 16055 15206 16069 15258
rect 16093 15206 16107 15258
rect 16107 15206 16119 15258
rect 16119 15206 16149 15258
rect 16173 15206 16183 15258
rect 16183 15206 16229 15258
rect 15933 15204 15989 15206
rect 16013 15204 16069 15206
rect 16093 15204 16149 15206
rect 16173 15204 16229 15206
rect 15273 14714 15329 14716
rect 15353 14714 15409 14716
rect 15433 14714 15489 14716
rect 15513 14714 15569 14716
rect 15273 14662 15319 14714
rect 15319 14662 15329 14714
rect 15353 14662 15383 14714
rect 15383 14662 15395 14714
rect 15395 14662 15409 14714
rect 15433 14662 15447 14714
rect 15447 14662 15459 14714
rect 15459 14662 15489 14714
rect 15513 14662 15523 14714
rect 15523 14662 15569 14714
rect 15273 14660 15329 14662
rect 15353 14660 15409 14662
rect 15433 14660 15489 14662
rect 15513 14660 15569 14662
rect 21000 20154 21056 20156
rect 21080 20154 21136 20156
rect 21160 20154 21216 20156
rect 21240 20154 21296 20156
rect 21000 20102 21046 20154
rect 21046 20102 21056 20154
rect 21080 20102 21110 20154
rect 21110 20102 21122 20154
rect 21122 20102 21136 20154
rect 21160 20102 21174 20154
rect 21174 20102 21186 20154
rect 21186 20102 21216 20154
rect 21240 20102 21250 20154
rect 21250 20102 21296 20154
rect 21000 20100 21056 20102
rect 21080 20100 21136 20102
rect 21160 20100 21216 20102
rect 21240 20100 21296 20102
rect 21660 19610 21716 19612
rect 21740 19610 21796 19612
rect 21820 19610 21876 19612
rect 21900 19610 21956 19612
rect 21660 19558 21706 19610
rect 21706 19558 21716 19610
rect 21740 19558 21770 19610
rect 21770 19558 21782 19610
rect 21782 19558 21796 19610
rect 21820 19558 21834 19610
rect 21834 19558 21846 19610
rect 21846 19558 21876 19610
rect 21900 19558 21910 19610
rect 21910 19558 21956 19610
rect 21660 19556 21716 19558
rect 21740 19556 21796 19558
rect 21820 19556 21876 19558
rect 21900 19556 21956 19558
rect 21000 19066 21056 19068
rect 21080 19066 21136 19068
rect 21160 19066 21216 19068
rect 21240 19066 21296 19068
rect 21000 19014 21046 19066
rect 21046 19014 21056 19066
rect 21080 19014 21110 19066
rect 21110 19014 21122 19066
rect 21122 19014 21136 19066
rect 21160 19014 21174 19066
rect 21174 19014 21186 19066
rect 21186 19014 21216 19066
rect 21240 19014 21250 19066
rect 21250 19014 21296 19066
rect 21000 19012 21056 19014
rect 21080 19012 21136 19014
rect 21160 19012 21216 19014
rect 21240 19012 21296 19014
rect 21660 18522 21716 18524
rect 21740 18522 21796 18524
rect 21820 18522 21876 18524
rect 21900 18522 21956 18524
rect 21660 18470 21706 18522
rect 21706 18470 21716 18522
rect 21740 18470 21770 18522
rect 21770 18470 21782 18522
rect 21782 18470 21796 18522
rect 21820 18470 21834 18522
rect 21834 18470 21846 18522
rect 21846 18470 21876 18522
rect 21900 18470 21910 18522
rect 21910 18470 21956 18522
rect 21660 18468 21716 18470
rect 21740 18468 21796 18470
rect 21820 18468 21876 18470
rect 21900 18468 21956 18470
rect 15933 14170 15989 14172
rect 16013 14170 16069 14172
rect 16093 14170 16149 14172
rect 16173 14170 16229 14172
rect 15933 14118 15979 14170
rect 15979 14118 15989 14170
rect 16013 14118 16043 14170
rect 16043 14118 16055 14170
rect 16055 14118 16069 14170
rect 16093 14118 16107 14170
rect 16107 14118 16119 14170
rect 16119 14118 16149 14170
rect 16173 14118 16183 14170
rect 16183 14118 16229 14170
rect 15933 14116 15989 14118
rect 16013 14116 16069 14118
rect 16093 14116 16149 14118
rect 16173 14116 16229 14118
rect 15273 13626 15329 13628
rect 15353 13626 15409 13628
rect 15433 13626 15489 13628
rect 15513 13626 15569 13628
rect 15273 13574 15319 13626
rect 15319 13574 15329 13626
rect 15353 13574 15383 13626
rect 15383 13574 15395 13626
rect 15395 13574 15409 13626
rect 15433 13574 15447 13626
rect 15447 13574 15459 13626
rect 15459 13574 15489 13626
rect 15513 13574 15523 13626
rect 15523 13574 15569 13626
rect 15273 13572 15329 13574
rect 15353 13572 15409 13574
rect 15433 13572 15489 13574
rect 15513 13572 15569 13574
rect 15273 12538 15329 12540
rect 15353 12538 15409 12540
rect 15433 12538 15489 12540
rect 15513 12538 15569 12540
rect 15273 12486 15319 12538
rect 15319 12486 15329 12538
rect 15353 12486 15383 12538
rect 15383 12486 15395 12538
rect 15395 12486 15409 12538
rect 15433 12486 15447 12538
rect 15447 12486 15459 12538
rect 15459 12486 15489 12538
rect 15513 12486 15523 12538
rect 15523 12486 15569 12538
rect 15273 12484 15329 12486
rect 15353 12484 15409 12486
rect 15433 12484 15489 12486
rect 15513 12484 15569 12486
rect 15273 11450 15329 11452
rect 15353 11450 15409 11452
rect 15433 11450 15489 11452
rect 15513 11450 15569 11452
rect 15273 11398 15319 11450
rect 15319 11398 15329 11450
rect 15353 11398 15383 11450
rect 15383 11398 15395 11450
rect 15395 11398 15409 11450
rect 15433 11398 15447 11450
rect 15447 11398 15459 11450
rect 15459 11398 15489 11450
rect 15513 11398 15523 11450
rect 15523 11398 15569 11450
rect 15273 11396 15329 11398
rect 15353 11396 15409 11398
rect 15433 11396 15489 11398
rect 15513 11396 15569 11398
rect 15933 13082 15989 13084
rect 16013 13082 16069 13084
rect 16093 13082 16149 13084
rect 16173 13082 16229 13084
rect 15933 13030 15979 13082
rect 15979 13030 15989 13082
rect 16013 13030 16043 13082
rect 16043 13030 16055 13082
rect 16055 13030 16069 13082
rect 16093 13030 16107 13082
rect 16107 13030 16119 13082
rect 16119 13030 16149 13082
rect 16173 13030 16183 13082
rect 16183 13030 16229 13082
rect 15933 13028 15989 13030
rect 16013 13028 16069 13030
rect 16093 13028 16149 13030
rect 16173 13028 16229 13030
rect 15933 11994 15989 11996
rect 16013 11994 16069 11996
rect 16093 11994 16149 11996
rect 16173 11994 16229 11996
rect 15933 11942 15979 11994
rect 15979 11942 15989 11994
rect 16013 11942 16043 11994
rect 16043 11942 16055 11994
rect 16055 11942 16069 11994
rect 16093 11942 16107 11994
rect 16107 11942 16119 11994
rect 16119 11942 16149 11994
rect 16173 11942 16183 11994
rect 16183 11942 16229 11994
rect 15933 11940 15989 11942
rect 16013 11940 16069 11942
rect 16093 11940 16149 11942
rect 16173 11940 16229 11942
rect 15933 10906 15989 10908
rect 16013 10906 16069 10908
rect 16093 10906 16149 10908
rect 16173 10906 16229 10908
rect 15933 10854 15979 10906
rect 15979 10854 15989 10906
rect 16013 10854 16043 10906
rect 16043 10854 16055 10906
rect 16055 10854 16069 10906
rect 16093 10854 16107 10906
rect 16107 10854 16119 10906
rect 16119 10854 16149 10906
rect 16173 10854 16183 10906
rect 16183 10854 16229 10906
rect 15933 10852 15989 10854
rect 16013 10852 16069 10854
rect 16093 10852 16149 10854
rect 16173 10852 16229 10854
rect 15273 10362 15329 10364
rect 15353 10362 15409 10364
rect 15433 10362 15489 10364
rect 15513 10362 15569 10364
rect 15273 10310 15319 10362
rect 15319 10310 15329 10362
rect 15353 10310 15383 10362
rect 15383 10310 15395 10362
rect 15395 10310 15409 10362
rect 15433 10310 15447 10362
rect 15447 10310 15459 10362
rect 15459 10310 15489 10362
rect 15513 10310 15523 10362
rect 15523 10310 15569 10362
rect 15273 10308 15329 10310
rect 15353 10308 15409 10310
rect 15433 10308 15489 10310
rect 15513 10308 15569 10310
rect 15273 9274 15329 9276
rect 15353 9274 15409 9276
rect 15433 9274 15489 9276
rect 15513 9274 15569 9276
rect 15273 9222 15319 9274
rect 15319 9222 15329 9274
rect 15353 9222 15383 9274
rect 15383 9222 15395 9274
rect 15395 9222 15409 9274
rect 15433 9222 15447 9274
rect 15447 9222 15459 9274
rect 15459 9222 15489 9274
rect 15513 9222 15523 9274
rect 15523 9222 15569 9274
rect 15273 9220 15329 9222
rect 15353 9220 15409 9222
rect 15433 9220 15489 9222
rect 15513 9220 15569 9222
rect 15273 8186 15329 8188
rect 15353 8186 15409 8188
rect 15433 8186 15489 8188
rect 15513 8186 15569 8188
rect 15273 8134 15319 8186
rect 15319 8134 15329 8186
rect 15353 8134 15383 8186
rect 15383 8134 15395 8186
rect 15395 8134 15409 8186
rect 15433 8134 15447 8186
rect 15447 8134 15459 8186
rect 15459 8134 15489 8186
rect 15513 8134 15523 8186
rect 15523 8134 15569 8186
rect 15273 8132 15329 8134
rect 15353 8132 15409 8134
rect 15433 8132 15489 8134
rect 15513 8132 15569 8134
rect 15933 9818 15989 9820
rect 16013 9818 16069 9820
rect 16093 9818 16149 9820
rect 16173 9818 16229 9820
rect 15933 9766 15979 9818
rect 15979 9766 15989 9818
rect 16013 9766 16043 9818
rect 16043 9766 16055 9818
rect 16055 9766 16069 9818
rect 16093 9766 16107 9818
rect 16107 9766 16119 9818
rect 16119 9766 16149 9818
rect 16173 9766 16183 9818
rect 16183 9766 16229 9818
rect 15933 9764 15989 9766
rect 16013 9764 16069 9766
rect 16093 9764 16149 9766
rect 16173 9764 16229 9766
rect 21000 17978 21056 17980
rect 21080 17978 21136 17980
rect 21160 17978 21216 17980
rect 21240 17978 21296 17980
rect 21000 17926 21046 17978
rect 21046 17926 21056 17978
rect 21080 17926 21110 17978
rect 21110 17926 21122 17978
rect 21122 17926 21136 17978
rect 21160 17926 21174 17978
rect 21174 17926 21186 17978
rect 21186 17926 21216 17978
rect 21240 17926 21250 17978
rect 21250 17926 21296 17978
rect 21000 17924 21056 17926
rect 21080 17924 21136 17926
rect 21160 17924 21216 17926
rect 21240 17924 21296 17926
rect 21660 17434 21716 17436
rect 21740 17434 21796 17436
rect 21820 17434 21876 17436
rect 21900 17434 21956 17436
rect 21660 17382 21706 17434
rect 21706 17382 21716 17434
rect 21740 17382 21770 17434
rect 21770 17382 21782 17434
rect 21782 17382 21796 17434
rect 21820 17382 21834 17434
rect 21834 17382 21846 17434
rect 21846 17382 21876 17434
rect 21900 17382 21910 17434
rect 21910 17382 21956 17434
rect 21660 17380 21716 17382
rect 21740 17380 21796 17382
rect 21820 17380 21876 17382
rect 21900 17380 21956 17382
rect 21000 16890 21056 16892
rect 21080 16890 21136 16892
rect 21160 16890 21216 16892
rect 21240 16890 21296 16892
rect 21000 16838 21046 16890
rect 21046 16838 21056 16890
rect 21080 16838 21110 16890
rect 21110 16838 21122 16890
rect 21122 16838 21136 16890
rect 21160 16838 21174 16890
rect 21174 16838 21186 16890
rect 21186 16838 21216 16890
rect 21240 16838 21250 16890
rect 21250 16838 21296 16890
rect 21000 16836 21056 16838
rect 21080 16836 21136 16838
rect 21160 16836 21216 16838
rect 21240 16836 21296 16838
rect 22006 16496 22062 16552
rect 21660 16346 21716 16348
rect 21740 16346 21796 16348
rect 21820 16346 21876 16348
rect 21900 16346 21956 16348
rect 21660 16294 21706 16346
rect 21706 16294 21716 16346
rect 21740 16294 21770 16346
rect 21770 16294 21782 16346
rect 21782 16294 21796 16346
rect 21820 16294 21834 16346
rect 21834 16294 21846 16346
rect 21846 16294 21876 16346
rect 21900 16294 21910 16346
rect 21910 16294 21956 16346
rect 21660 16292 21716 16294
rect 21740 16292 21796 16294
rect 21820 16292 21876 16294
rect 21900 16292 21956 16294
rect 23662 22480 23718 22536
rect 23386 20440 23442 20496
rect 21000 15802 21056 15804
rect 21080 15802 21136 15804
rect 21160 15802 21216 15804
rect 21240 15802 21296 15804
rect 21000 15750 21046 15802
rect 21046 15750 21056 15802
rect 21080 15750 21110 15802
rect 21110 15750 21122 15802
rect 21122 15750 21136 15802
rect 21160 15750 21174 15802
rect 21174 15750 21186 15802
rect 21186 15750 21216 15802
rect 21240 15750 21250 15802
rect 21250 15750 21296 15802
rect 21000 15748 21056 15750
rect 21080 15748 21136 15750
rect 21160 15748 21216 15750
rect 21240 15748 21296 15750
rect 21000 14714 21056 14716
rect 21080 14714 21136 14716
rect 21160 14714 21216 14716
rect 21240 14714 21296 14716
rect 21000 14662 21046 14714
rect 21046 14662 21056 14714
rect 21080 14662 21110 14714
rect 21110 14662 21122 14714
rect 21122 14662 21136 14714
rect 21160 14662 21174 14714
rect 21174 14662 21186 14714
rect 21186 14662 21216 14714
rect 21240 14662 21250 14714
rect 21250 14662 21296 14714
rect 21000 14660 21056 14662
rect 21080 14660 21136 14662
rect 21160 14660 21216 14662
rect 21240 14660 21296 14662
rect 21660 15258 21716 15260
rect 21740 15258 21796 15260
rect 21820 15258 21876 15260
rect 21900 15258 21956 15260
rect 21660 15206 21706 15258
rect 21706 15206 21716 15258
rect 21740 15206 21770 15258
rect 21770 15206 21782 15258
rect 21782 15206 21796 15258
rect 21820 15206 21834 15258
rect 21834 15206 21846 15258
rect 21846 15206 21876 15258
rect 21900 15206 21910 15258
rect 21910 15206 21956 15258
rect 21660 15204 21716 15206
rect 21740 15204 21796 15206
rect 21820 15204 21876 15206
rect 21900 15204 21956 15206
rect 23386 19080 23442 19136
rect 23294 18400 23350 18456
rect 23662 21800 23718 21856
rect 23662 21120 23718 21176
rect 23662 19760 23718 19816
rect 23662 17756 23664 17776
rect 23664 17756 23716 17776
rect 23716 17756 23718 17776
rect 23662 17720 23718 17756
rect 23662 17060 23718 17096
rect 23662 17040 23664 17060
rect 23664 17040 23716 17060
rect 23716 17040 23718 17060
rect 23202 16496 23258 16552
rect 23386 15000 23442 15056
rect 21660 14170 21716 14172
rect 21740 14170 21796 14172
rect 21820 14170 21876 14172
rect 21900 14170 21956 14172
rect 21660 14118 21706 14170
rect 21706 14118 21716 14170
rect 21740 14118 21770 14170
rect 21770 14118 21782 14170
rect 21782 14118 21796 14170
rect 21820 14118 21834 14170
rect 21834 14118 21846 14170
rect 21846 14118 21876 14170
rect 21900 14118 21910 14170
rect 21910 14118 21956 14170
rect 21660 14116 21716 14118
rect 21740 14116 21796 14118
rect 21820 14116 21876 14118
rect 21900 14116 21956 14118
rect 21000 13626 21056 13628
rect 21080 13626 21136 13628
rect 21160 13626 21216 13628
rect 21240 13626 21296 13628
rect 21000 13574 21046 13626
rect 21046 13574 21056 13626
rect 21080 13574 21110 13626
rect 21110 13574 21122 13626
rect 21122 13574 21136 13626
rect 21160 13574 21174 13626
rect 21174 13574 21186 13626
rect 21186 13574 21216 13626
rect 21240 13574 21250 13626
rect 21250 13574 21296 13626
rect 21000 13572 21056 13574
rect 21080 13572 21136 13574
rect 21160 13572 21216 13574
rect 21240 13572 21296 13574
rect 21660 13082 21716 13084
rect 21740 13082 21796 13084
rect 21820 13082 21876 13084
rect 21900 13082 21956 13084
rect 21660 13030 21706 13082
rect 21706 13030 21716 13082
rect 21740 13030 21770 13082
rect 21770 13030 21782 13082
rect 21782 13030 21796 13082
rect 21820 13030 21834 13082
rect 21834 13030 21846 13082
rect 21846 13030 21876 13082
rect 21900 13030 21910 13082
rect 21910 13030 21956 13082
rect 21660 13028 21716 13030
rect 21740 13028 21796 13030
rect 21820 13028 21876 13030
rect 21900 13028 21956 13030
rect 21000 12538 21056 12540
rect 21080 12538 21136 12540
rect 21160 12538 21216 12540
rect 21240 12538 21296 12540
rect 21000 12486 21046 12538
rect 21046 12486 21056 12538
rect 21080 12486 21110 12538
rect 21110 12486 21122 12538
rect 21122 12486 21136 12538
rect 21160 12486 21174 12538
rect 21174 12486 21186 12538
rect 21186 12486 21216 12538
rect 21240 12486 21250 12538
rect 21250 12486 21296 12538
rect 21000 12484 21056 12486
rect 21080 12484 21136 12486
rect 21160 12484 21216 12486
rect 21240 12484 21296 12486
rect 23662 16360 23718 16416
rect 23662 15680 23718 15736
rect 23662 14320 23718 14376
rect 23386 13640 23442 13696
rect 23662 12960 23718 13016
rect 21660 11994 21716 11996
rect 21740 11994 21796 11996
rect 21820 11994 21876 11996
rect 21900 11994 21956 11996
rect 21660 11942 21706 11994
rect 21706 11942 21716 11994
rect 21740 11942 21770 11994
rect 21770 11942 21782 11994
rect 21782 11942 21796 11994
rect 21820 11942 21834 11994
rect 21834 11942 21846 11994
rect 21846 11942 21876 11994
rect 21900 11942 21910 11994
rect 21910 11942 21956 11994
rect 21660 11940 21716 11942
rect 21740 11940 21796 11942
rect 21820 11940 21876 11942
rect 21900 11940 21956 11942
rect 15933 8730 15989 8732
rect 16013 8730 16069 8732
rect 16093 8730 16149 8732
rect 16173 8730 16229 8732
rect 15933 8678 15979 8730
rect 15979 8678 15989 8730
rect 16013 8678 16043 8730
rect 16043 8678 16055 8730
rect 16055 8678 16069 8730
rect 16093 8678 16107 8730
rect 16107 8678 16119 8730
rect 16119 8678 16149 8730
rect 16173 8678 16183 8730
rect 16183 8678 16229 8730
rect 15933 8676 15989 8678
rect 16013 8676 16069 8678
rect 16093 8676 16149 8678
rect 16173 8676 16229 8678
rect 15933 7642 15989 7644
rect 16013 7642 16069 7644
rect 16093 7642 16149 7644
rect 16173 7642 16229 7644
rect 15933 7590 15979 7642
rect 15979 7590 15989 7642
rect 16013 7590 16043 7642
rect 16043 7590 16055 7642
rect 16055 7590 16069 7642
rect 16093 7590 16107 7642
rect 16107 7590 16119 7642
rect 16119 7590 16149 7642
rect 16173 7590 16183 7642
rect 16183 7590 16229 7642
rect 15933 7588 15989 7590
rect 16013 7588 16069 7590
rect 16093 7588 16149 7590
rect 16173 7588 16229 7590
rect 15273 7098 15329 7100
rect 15353 7098 15409 7100
rect 15433 7098 15489 7100
rect 15513 7098 15569 7100
rect 15273 7046 15319 7098
rect 15319 7046 15329 7098
rect 15353 7046 15383 7098
rect 15383 7046 15395 7098
rect 15395 7046 15409 7098
rect 15433 7046 15447 7098
rect 15447 7046 15459 7098
rect 15459 7046 15489 7098
rect 15513 7046 15523 7098
rect 15523 7046 15569 7098
rect 15273 7044 15329 7046
rect 15353 7044 15409 7046
rect 15433 7044 15489 7046
rect 15513 7044 15569 7046
rect 15273 6010 15329 6012
rect 15353 6010 15409 6012
rect 15433 6010 15489 6012
rect 15513 6010 15569 6012
rect 15273 5958 15319 6010
rect 15319 5958 15329 6010
rect 15353 5958 15383 6010
rect 15383 5958 15395 6010
rect 15395 5958 15409 6010
rect 15433 5958 15447 6010
rect 15447 5958 15459 6010
rect 15459 5958 15489 6010
rect 15513 5958 15523 6010
rect 15523 5958 15569 6010
rect 15273 5956 15329 5958
rect 15353 5956 15409 5958
rect 15433 5956 15489 5958
rect 15513 5956 15569 5958
rect 15273 4922 15329 4924
rect 15353 4922 15409 4924
rect 15433 4922 15489 4924
rect 15513 4922 15569 4924
rect 15273 4870 15319 4922
rect 15319 4870 15329 4922
rect 15353 4870 15383 4922
rect 15383 4870 15395 4922
rect 15395 4870 15409 4922
rect 15433 4870 15447 4922
rect 15447 4870 15459 4922
rect 15459 4870 15489 4922
rect 15513 4870 15523 4922
rect 15523 4870 15569 4922
rect 15273 4868 15329 4870
rect 15353 4868 15409 4870
rect 15433 4868 15489 4870
rect 15513 4868 15569 4870
rect 15933 6554 15989 6556
rect 16013 6554 16069 6556
rect 16093 6554 16149 6556
rect 16173 6554 16229 6556
rect 15933 6502 15979 6554
rect 15979 6502 15989 6554
rect 16013 6502 16043 6554
rect 16043 6502 16055 6554
rect 16055 6502 16069 6554
rect 16093 6502 16107 6554
rect 16107 6502 16119 6554
rect 16119 6502 16149 6554
rect 16173 6502 16183 6554
rect 16183 6502 16229 6554
rect 15933 6500 15989 6502
rect 16013 6500 16069 6502
rect 16093 6500 16149 6502
rect 16173 6500 16229 6502
rect 15933 5466 15989 5468
rect 16013 5466 16069 5468
rect 16093 5466 16149 5468
rect 16173 5466 16229 5468
rect 15933 5414 15979 5466
rect 15979 5414 15989 5466
rect 16013 5414 16043 5466
rect 16043 5414 16055 5466
rect 16055 5414 16069 5466
rect 16093 5414 16107 5466
rect 16107 5414 16119 5466
rect 16119 5414 16149 5466
rect 16173 5414 16183 5466
rect 16183 5414 16229 5466
rect 15933 5412 15989 5414
rect 16013 5412 16069 5414
rect 16093 5412 16149 5414
rect 16173 5412 16229 5414
rect 15933 4378 15989 4380
rect 16013 4378 16069 4380
rect 16093 4378 16149 4380
rect 16173 4378 16229 4380
rect 15933 4326 15979 4378
rect 15979 4326 15989 4378
rect 16013 4326 16043 4378
rect 16043 4326 16055 4378
rect 16055 4326 16069 4378
rect 16093 4326 16107 4378
rect 16107 4326 16119 4378
rect 16119 4326 16149 4378
rect 16173 4326 16183 4378
rect 16183 4326 16229 4378
rect 15933 4324 15989 4326
rect 16013 4324 16069 4326
rect 16093 4324 16149 4326
rect 16173 4324 16229 4326
rect 15273 3834 15329 3836
rect 15353 3834 15409 3836
rect 15433 3834 15489 3836
rect 15513 3834 15569 3836
rect 15273 3782 15319 3834
rect 15319 3782 15329 3834
rect 15353 3782 15383 3834
rect 15383 3782 15395 3834
rect 15395 3782 15409 3834
rect 15433 3782 15447 3834
rect 15447 3782 15459 3834
rect 15459 3782 15489 3834
rect 15513 3782 15523 3834
rect 15523 3782 15569 3834
rect 15273 3780 15329 3782
rect 15353 3780 15409 3782
rect 15433 3780 15489 3782
rect 15513 3780 15569 3782
rect 15273 2746 15329 2748
rect 15353 2746 15409 2748
rect 15433 2746 15489 2748
rect 15513 2746 15569 2748
rect 15273 2694 15319 2746
rect 15319 2694 15329 2746
rect 15353 2694 15383 2746
rect 15383 2694 15395 2746
rect 15395 2694 15409 2746
rect 15433 2694 15447 2746
rect 15447 2694 15459 2746
rect 15459 2694 15489 2746
rect 15513 2694 15523 2746
rect 15523 2694 15569 2746
rect 15273 2692 15329 2694
rect 15353 2692 15409 2694
rect 15433 2692 15489 2694
rect 15513 2692 15569 2694
rect 15933 3290 15989 3292
rect 16013 3290 16069 3292
rect 16093 3290 16149 3292
rect 16173 3290 16229 3292
rect 15933 3238 15979 3290
rect 15979 3238 15989 3290
rect 16013 3238 16043 3290
rect 16043 3238 16055 3290
rect 16055 3238 16069 3290
rect 16093 3238 16107 3290
rect 16107 3238 16119 3290
rect 16119 3238 16149 3290
rect 16173 3238 16183 3290
rect 16183 3238 16229 3290
rect 15933 3236 15989 3238
rect 16013 3236 16069 3238
rect 16093 3236 16149 3238
rect 16173 3236 16229 3238
rect 21000 11450 21056 11452
rect 21080 11450 21136 11452
rect 21160 11450 21216 11452
rect 21240 11450 21296 11452
rect 21000 11398 21046 11450
rect 21046 11398 21056 11450
rect 21080 11398 21110 11450
rect 21110 11398 21122 11450
rect 21122 11398 21136 11450
rect 21160 11398 21174 11450
rect 21174 11398 21186 11450
rect 21186 11398 21216 11450
rect 21240 11398 21250 11450
rect 21250 11398 21296 11450
rect 21000 11396 21056 11398
rect 21080 11396 21136 11398
rect 21160 11396 21216 11398
rect 21240 11396 21296 11398
rect 21000 10362 21056 10364
rect 21080 10362 21136 10364
rect 21160 10362 21216 10364
rect 21240 10362 21296 10364
rect 21000 10310 21046 10362
rect 21046 10310 21056 10362
rect 21080 10310 21110 10362
rect 21110 10310 21122 10362
rect 21122 10310 21136 10362
rect 21160 10310 21174 10362
rect 21174 10310 21186 10362
rect 21186 10310 21216 10362
rect 21240 10310 21250 10362
rect 21250 10310 21296 10362
rect 21000 10308 21056 10310
rect 21080 10308 21136 10310
rect 21160 10308 21216 10310
rect 21240 10308 21296 10310
rect 21000 9274 21056 9276
rect 21080 9274 21136 9276
rect 21160 9274 21216 9276
rect 21240 9274 21296 9276
rect 21000 9222 21046 9274
rect 21046 9222 21056 9274
rect 21080 9222 21110 9274
rect 21110 9222 21122 9274
rect 21122 9222 21136 9274
rect 21160 9222 21174 9274
rect 21174 9222 21186 9274
rect 21186 9222 21216 9274
rect 21240 9222 21250 9274
rect 21250 9222 21296 9274
rect 21000 9220 21056 9222
rect 21080 9220 21136 9222
rect 21160 9220 21216 9222
rect 21240 9220 21296 9222
rect 21000 8186 21056 8188
rect 21080 8186 21136 8188
rect 21160 8186 21216 8188
rect 21240 8186 21296 8188
rect 21000 8134 21046 8186
rect 21046 8134 21056 8186
rect 21080 8134 21110 8186
rect 21110 8134 21122 8186
rect 21122 8134 21136 8186
rect 21160 8134 21174 8186
rect 21174 8134 21186 8186
rect 21186 8134 21216 8186
rect 21240 8134 21250 8186
rect 21250 8134 21296 8186
rect 21000 8132 21056 8134
rect 21080 8132 21136 8134
rect 21160 8132 21216 8134
rect 21240 8132 21296 8134
rect 21660 10906 21716 10908
rect 21740 10906 21796 10908
rect 21820 10906 21876 10908
rect 21900 10906 21956 10908
rect 21660 10854 21706 10906
rect 21706 10854 21716 10906
rect 21740 10854 21770 10906
rect 21770 10854 21782 10906
rect 21782 10854 21796 10906
rect 21820 10854 21834 10906
rect 21834 10854 21846 10906
rect 21846 10854 21876 10906
rect 21900 10854 21910 10906
rect 21910 10854 21956 10906
rect 21660 10852 21716 10854
rect 21740 10852 21796 10854
rect 21820 10852 21876 10854
rect 21900 10852 21956 10854
rect 23386 12280 23442 12336
rect 23662 11600 23718 11656
rect 21660 9818 21716 9820
rect 21740 9818 21796 9820
rect 21820 9818 21876 9820
rect 21900 9818 21956 9820
rect 21660 9766 21706 9818
rect 21706 9766 21716 9818
rect 21740 9766 21770 9818
rect 21770 9766 21782 9818
rect 21782 9766 21796 9818
rect 21820 9766 21834 9818
rect 21834 9766 21846 9818
rect 21846 9766 21876 9818
rect 21900 9766 21910 9818
rect 21910 9766 21956 9818
rect 21660 9764 21716 9766
rect 21740 9764 21796 9766
rect 21820 9764 21876 9766
rect 21900 9764 21956 9766
rect 21660 8730 21716 8732
rect 21740 8730 21796 8732
rect 21820 8730 21876 8732
rect 21900 8730 21956 8732
rect 21660 8678 21706 8730
rect 21706 8678 21716 8730
rect 21740 8678 21770 8730
rect 21770 8678 21782 8730
rect 21782 8678 21796 8730
rect 21820 8678 21834 8730
rect 21834 8678 21846 8730
rect 21846 8678 21876 8730
rect 21900 8678 21910 8730
rect 21910 8678 21956 8730
rect 21660 8676 21716 8678
rect 21740 8676 21796 8678
rect 21820 8676 21876 8678
rect 21900 8676 21956 8678
rect 21000 7098 21056 7100
rect 21080 7098 21136 7100
rect 21160 7098 21216 7100
rect 21240 7098 21296 7100
rect 21000 7046 21046 7098
rect 21046 7046 21056 7098
rect 21080 7046 21110 7098
rect 21110 7046 21122 7098
rect 21122 7046 21136 7098
rect 21160 7046 21174 7098
rect 21174 7046 21186 7098
rect 21186 7046 21216 7098
rect 21240 7046 21250 7098
rect 21250 7046 21296 7098
rect 21000 7044 21056 7046
rect 21080 7044 21136 7046
rect 21160 7044 21216 7046
rect 21240 7044 21296 7046
rect 21660 7642 21716 7644
rect 21740 7642 21796 7644
rect 21820 7642 21876 7644
rect 21900 7642 21956 7644
rect 21660 7590 21706 7642
rect 21706 7590 21716 7642
rect 21740 7590 21770 7642
rect 21770 7590 21782 7642
rect 21782 7590 21796 7642
rect 21820 7590 21834 7642
rect 21834 7590 21846 7642
rect 21846 7590 21876 7642
rect 21900 7590 21910 7642
rect 21910 7590 21956 7642
rect 21660 7588 21716 7590
rect 21740 7588 21796 7590
rect 21820 7588 21876 7590
rect 21900 7588 21956 7590
rect 21000 6010 21056 6012
rect 21080 6010 21136 6012
rect 21160 6010 21216 6012
rect 21240 6010 21296 6012
rect 21000 5958 21046 6010
rect 21046 5958 21056 6010
rect 21080 5958 21110 6010
rect 21110 5958 21122 6010
rect 21122 5958 21136 6010
rect 21160 5958 21174 6010
rect 21174 5958 21186 6010
rect 21186 5958 21216 6010
rect 21240 5958 21250 6010
rect 21250 5958 21296 6010
rect 21000 5956 21056 5958
rect 21080 5956 21136 5958
rect 21160 5956 21216 5958
rect 21240 5956 21296 5958
rect 21000 4922 21056 4924
rect 21080 4922 21136 4924
rect 21160 4922 21216 4924
rect 21240 4922 21296 4924
rect 21000 4870 21046 4922
rect 21046 4870 21056 4922
rect 21080 4870 21110 4922
rect 21110 4870 21122 4922
rect 21122 4870 21136 4922
rect 21160 4870 21174 4922
rect 21174 4870 21186 4922
rect 21186 4870 21216 4922
rect 21240 4870 21250 4922
rect 21250 4870 21296 4922
rect 21000 4868 21056 4870
rect 21080 4868 21136 4870
rect 21160 4868 21216 4870
rect 21240 4868 21296 4870
rect 21000 3834 21056 3836
rect 21080 3834 21136 3836
rect 21160 3834 21216 3836
rect 21240 3834 21296 3836
rect 21000 3782 21046 3834
rect 21046 3782 21056 3834
rect 21080 3782 21110 3834
rect 21110 3782 21122 3834
rect 21122 3782 21136 3834
rect 21160 3782 21174 3834
rect 21174 3782 21186 3834
rect 21186 3782 21216 3834
rect 21240 3782 21250 3834
rect 21250 3782 21296 3834
rect 21000 3780 21056 3782
rect 21080 3780 21136 3782
rect 21160 3780 21216 3782
rect 21240 3780 21296 3782
rect 21660 6554 21716 6556
rect 21740 6554 21796 6556
rect 21820 6554 21876 6556
rect 21900 6554 21956 6556
rect 21660 6502 21706 6554
rect 21706 6502 21716 6554
rect 21740 6502 21770 6554
rect 21770 6502 21782 6554
rect 21782 6502 21796 6554
rect 21820 6502 21834 6554
rect 21834 6502 21846 6554
rect 21846 6502 21876 6554
rect 21900 6502 21910 6554
rect 21910 6502 21956 6554
rect 21660 6500 21716 6502
rect 21740 6500 21796 6502
rect 21820 6500 21876 6502
rect 21900 6500 21956 6502
rect 21660 5466 21716 5468
rect 21740 5466 21796 5468
rect 21820 5466 21876 5468
rect 21900 5466 21956 5468
rect 21660 5414 21706 5466
rect 21706 5414 21716 5466
rect 21740 5414 21770 5466
rect 21770 5414 21782 5466
rect 21782 5414 21796 5466
rect 21820 5414 21834 5466
rect 21834 5414 21846 5466
rect 21846 5414 21876 5466
rect 21900 5414 21910 5466
rect 21910 5414 21956 5466
rect 21660 5412 21716 5414
rect 21740 5412 21796 5414
rect 21820 5412 21876 5414
rect 21900 5412 21956 5414
rect 23386 10920 23442 10976
rect 23662 10240 23718 10296
rect 23386 8200 23442 8256
rect 23662 9560 23718 9616
rect 23662 8880 23718 8936
rect 23662 7520 23718 7576
rect 23662 6840 23718 6896
rect 23662 6160 23718 6216
rect 23386 5480 23442 5536
rect 23662 4800 23718 4856
rect 21660 4378 21716 4380
rect 21740 4378 21796 4380
rect 21820 4378 21876 4380
rect 21900 4378 21956 4380
rect 21660 4326 21706 4378
rect 21706 4326 21716 4378
rect 21740 4326 21770 4378
rect 21770 4326 21782 4378
rect 21782 4326 21796 4378
rect 21820 4326 21834 4378
rect 21834 4326 21846 4378
rect 21846 4326 21876 4378
rect 21900 4326 21910 4378
rect 21910 4326 21956 4378
rect 21660 4324 21716 4326
rect 21740 4324 21796 4326
rect 21820 4324 21876 4326
rect 21900 4324 21956 4326
rect 21660 3290 21716 3292
rect 21740 3290 21796 3292
rect 21820 3290 21876 3292
rect 21900 3290 21956 3292
rect 21660 3238 21706 3290
rect 21706 3238 21716 3290
rect 21740 3238 21770 3290
rect 21770 3238 21782 3290
rect 21782 3238 21796 3290
rect 21820 3238 21834 3290
rect 21834 3238 21846 3290
rect 21846 3238 21876 3290
rect 21900 3238 21910 3290
rect 21910 3238 21956 3290
rect 21660 3236 21716 3238
rect 21740 3236 21796 3238
rect 21820 3236 21876 3238
rect 21900 3236 21956 3238
rect 23662 4120 23718 4176
rect 23662 3476 23664 3496
rect 23664 3476 23716 3496
rect 23716 3476 23718 3496
rect 23662 3440 23718 3476
rect 23662 2760 23718 2816
rect 21000 2746 21056 2748
rect 21080 2746 21136 2748
rect 21160 2746 21216 2748
rect 21240 2746 21296 2748
rect 21000 2694 21046 2746
rect 21046 2694 21056 2746
rect 21080 2694 21110 2746
rect 21110 2694 21122 2746
rect 21122 2694 21136 2746
rect 21160 2694 21174 2746
rect 21174 2694 21186 2746
rect 21186 2694 21216 2746
rect 21240 2694 21250 2746
rect 21250 2694 21296 2746
rect 21000 2692 21056 2694
rect 21080 2692 21136 2694
rect 21160 2692 21216 2694
rect 21240 2692 21296 2694
rect 15933 2202 15989 2204
rect 16013 2202 16069 2204
rect 16093 2202 16149 2204
rect 16173 2202 16229 2204
rect 15933 2150 15979 2202
rect 15979 2150 15989 2202
rect 16013 2150 16043 2202
rect 16043 2150 16055 2202
rect 16055 2150 16069 2202
rect 16093 2150 16107 2202
rect 16107 2150 16119 2202
rect 16119 2150 16149 2202
rect 16173 2150 16183 2202
rect 16183 2150 16229 2202
rect 15933 2148 15989 2150
rect 16013 2148 16069 2150
rect 16093 2148 16149 2150
rect 16173 2148 16229 2150
rect 21660 2202 21716 2204
rect 21740 2202 21796 2204
rect 21820 2202 21876 2204
rect 21900 2202 21956 2204
rect 21660 2150 21706 2202
rect 21706 2150 21716 2202
rect 21740 2150 21770 2202
rect 21770 2150 21782 2202
rect 21782 2150 21796 2202
rect 21820 2150 21834 2202
rect 21834 2150 21846 2202
rect 21846 2150 21876 2202
rect 21900 2150 21910 2202
rect 21910 2150 21956 2202
rect 21660 2148 21716 2150
rect 21740 2148 21796 2150
rect 21820 2148 21876 2150
rect 21900 2148 21956 2150
<< metal3 >>
rect 4469 25056 4785 25057
rect 4469 24992 4475 25056
rect 4539 24992 4555 25056
rect 4619 24992 4635 25056
rect 4699 24992 4715 25056
rect 4779 24992 4785 25056
rect 4469 24991 4785 24992
rect 10196 25056 10512 25057
rect 10196 24992 10202 25056
rect 10266 24992 10282 25056
rect 10346 24992 10362 25056
rect 10426 24992 10442 25056
rect 10506 24992 10512 25056
rect 10196 24991 10512 24992
rect 15923 25056 16239 25057
rect 15923 24992 15929 25056
rect 15993 24992 16009 25056
rect 16073 24992 16089 25056
rect 16153 24992 16169 25056
rect 16233 24992 16239 25056
rect 15923 24991 16239 24992
rect 21650 25056 21966 25057
rect 21650 24992 21656 25056
rect 21720 24992 21736 25056
rect 21800 24992 21816 25056
rect 21880 24992 21896 25056
rect 21960 24992 21966 25056
rect 21650 24991 21966 24992
rect 23657 24578 23723 24581
rect 24372 24578 25172 24608
rect 23657 24576 25172 24578
rect 23657 24520 23662 24576
rect 23718 24520 25172 24576
rect 23657 24518 25172 24520
rect 23657 24515 23723 24518
rect 3809 24512 4125 24513
rect 3809 24448 3815 24512
rect 3879 24448 3895 24512
rect 3959 24448 3975 24512
rect 4039 24448 4055 24512
rect 4119 24448 4125 24512
rect 3809 24447 4125 24448
rect 9536 24512 9852 24513
rect 9536 24448 9542 24512
rect 9606 24448 9622 24512
rect 9686 24448 9702 24512
rect 9766 24448 9782 24512
rect 9846 24448 9852 24512
rect 9536 24447 9852 24448
rect 15263 24512 15579 24513
rect 15263 24448 15269 24512
rect 15333 24448 15349 24512
rect 15413 24448 15429 24512
rect 15493 24448 15509 24512
rect 15573 24448 15579 24512
rect 15263 24447 15579 24448
rect 20990 24512 21306 24513
rect 20990 24448 20996 24512
rect 21060 24448 21076 24512
rect 21140 24448 21156 24512
rect 21220 24448 21236 24512
rect 21300 24448 21306 24512
rect 24372 24488 25172 24518
rect 20990 24447 21306 24448
rect 4469 23968 4785 23969
rect 4469 23904 4475 23968
rect 4539 23904 4555 23968
rect 4619 23904 4635 23968
rect 4699 23904 4715 23968
rect 4779 23904 4785 23968
rect 4469 23903 4785 23904
rect 10196 23968 10512 23969
rect 10196 23904 10202 23968
rect 10266 23904 10282 23968
rect 10346 23904 10362 23968
rect 10426 23904 10442 23968
rect 10506 23904 10512 23968
rect 10196 23903 10512 23904
rect 15923 23968 16239 23969
rect 15923 23904 15929 23968
rect 15993 23904 16009 23968
rect 16073 23904 16089 23968
rect 16153 23904 16169 23968
rect 16233 23904 16239 23968
rect 15923 23903 16239 23904
rect 21650 23968 21966 23969
rect 21650 23904 21656 23968
rect 21720 23904 21736 23968
rect 21800 23904 21816 23968
rect 21880 23904 21896 23968
rect 21960 23904 21966 23968
rect 21650 23903 21966 23904
rect 23657 23898 23723 23901
rect 24372 23898 25172 23928
rect 23657 23896 25172 23898
rect 23657 23840 23662 23896
rect 23718 23840 25172 23896
rect 23657 23838 25172 23840
rect 23657 23835 23723 23838
rect 24372 23808 25172 23838
rect 3809 23424 4125 23425
rect 3809 23360 3815 23424
rect 3879 23360 3895 23424
rect 3959 23360 3975 23424
rect 4039 23360 4055 23424
rect 4119 23360 4125 23424
rect 3809 23359 4125 23360
rect 9536 23424 9852 23425
rect 9536 23360 9542 23424
rect 9606 23360 9622 23424
rect 9686 23360 9702 23424
rect 9766 23360 9782 23424
rect 9846 23360 9852 23424
rect 9536 23359 9852 23360
rect 15263 23424 15579 23425
rect 15263 23360 15269 23424
rect 15333 23360 15349 23424
rect 15413 23360 15429 23424
rect 15493 23360 15509 23424
rect 15573 23360 15579 23424
rect 15263 23359 15579 23360
rect 20990 23424 21306 23425
rect 20990 23360 20996 23424
rect 21060 23360 21076 23424
rect 21140 23360 21156 23424
rect 21220 23360 21236 23424
rect 21300 23360 21306 23424
rect 20990 23359 21306 23360
rect 23381 23218 23447 23221
rect 24372 23218 25172 23248
rect 23381 23216 25172 23218
rect 23381 23160 23386 23216
rect 23442 23160 25172 23216
rect 23381 23158 25172 23160
rect 23381 23155 23447 23158
rect 24372 23128 25172 23158
rect 4469 22880 4785 22881
rect 4469 22816 4475 22880
rect 4539 22816 4555 22880
rect 4619 22816 4635 22880
rect 4699 22816 4715 22880
rect 4779 22816 4785 22880
rect 4469 22815 4785 22816
rect 10196 22880 10512 22881
rect 10196 22816 10202 22880
rect 10266 22816 10282 22880
rect 10346 22816 10362 22880
rect 10426 22816 10442 22880
rect 10506 22816 10512 22880
rect 10196 22815 10512 22816
rect 15923 22880 16239 22881
rect 15923 22816 15929 22880
rect 15993 22816 16009 22880
rect 16073 22816 16089 22880
rect 16153 22816 16169 22880
rect 16233 22816 16239 22880
rect 15923 22815 16239 22816
rect 21650 22880 21966 22881
rect 21650 22816 21656 22880
rect 21720 22816 21736 22880
rect 21800 22816 21816 22880
rect 21880 22816 21896 22880
rect 21960 22816 21966 22880
rect 21650 22815 21966 22816
rect 23657 22538 23723 22541
rect 24372 22538 25172 22568
rect 23657 22536 25172 22538
rect 23657 22480 23662 22536
rect 23718 22480 25172 22536
rect 23657 22478 25172 22480
rect 23657 22475 23723 22478
rect 24372 22448 25172 22478
rect 3809 22336 4125 22337
rect 3809 22272 3815 22336
rect 3879 22272 3895 22336
rect 3959 22272 3975 22336
rect 4039 22272 4055 22336
rect 4119 22272 4125 22336
rect 3809 22271 4125 22272
rect 9536 22336 9852 22337
rect 9536 22272 9542 22336
rect 9606 22272 9622 22336
rect 9686 22272 9702 22336
rect 9766 22272 9782 22336
rect 9846 22272 9852 22336
rect 9536 22271 9852 22272
rect 15263 22336 15579 22337
rect 15263 22272 15269 22336
rect 15333 22272 15349 22336
rect 15413 22272 15429 22336
rect 15493 22272 15509 22336
rect 15573 22272 15579 22336
rect 15263 22271 15579 22272
rect 20990 22336 21306 22337
rect 20990 22272 20996 22336
rect 21060 22272 21076 22336
rect 21140 22272 21156 22336
rect 21220 22272 21236 22336
rect 21300 22272 21306 22336
rect 20990 22271 21306 22272
rect 23657 21858 23723 21861
rect 24372 21858 25172 21888
rect 23657 21856 25172 21858
rect 23657 21800 23662 21856
rect 23718 21800 25172 21856
rect 23657 21798 25172 21800
rect 23657 21795 23723 21798
rect 4469 21792 4785 21793
rect 4469 21728 4475 21792
rect 4539 21728 4555 21792
rect 4619 21728 4635 21792
rect 4699 21728 4715 21792
rect 4779 21728 4785 21792
rect 4469 21727 4785 21728
rect 10196 21792 10512 21793
rect 10196 21728 10202 21792
rect 10266 21728 10282 21792
rect 10346 21728 10362 21792
rect 10426 21728 10442 21792
rect 10506 21728 10512 21792
rect 10196 21727 10512 21728
rect 15923 21792 16239 21793
rect 15923 21728 15929 21792
rect 15993 21728 16009 21792
rect 16073 21728 16089 21792
rect 16153 21728 16169 21792
rect 16233 21728 16239 21792
rect 15923 21727 16239 21728
rect 21650 21792 21966 21793
rect 21650 21728 21656 21792
rect 21720 21728 21736 21792
rect 21800 21728 21816 21792
rect 21880 21728 21896 21792
rect 21960 21728 21966 21792
rect 24372 21768 25172 21798
rect 21650 21727 21966 21728
rect 841 21314 907 21317
rect 798 21312 907 21314
rect 798 21256 846 21312
rect 902 21256 907 21312
rect 798 21251 907 21256
rect 798 21208 858 21251
rect 0 21118 858 21208
rect 3809 21248 4125 21249
rect 3809 21184 3815 21248
rect 3879 21184 3895 21248
rect 3959 21184 3975 21248
rect 4039 21184 4055 21248
rect 4119 21184 4125 21248
rect 3809 21183 4125 21184
rect 9536 21248 9852 21249
rect 9536 21184 9542 21248
rect 9606 21184 9622 21248
rect 9686 21184 9702 21248
rect 9766 21184 9782 21248
rect 9846 21184 9852 21248
rect 9536 21183 9852 21184
rect 15263 21248 15579 21249
rect 15263 21184 15269 21248
rect 15333 21184 15349 21248
rect 15413 21184 15429 21248
rect 15493 21184 15509 21248
rect 15573 21184 15579 21248
rect 15263 21183 15579 21184
rect 20990 21248 21306 21249
rect 20990 21184 20996 21248
rect 21060 21184 21076 21248
rect 21140 21184 21156 21248
rect 21220 21184 21236 21248
rect 21300 21184 21306 21248
rect 20990 21183 21306 21184
rect 23657 21178 23723 21181
rect 24372 21178 25172 21208
rect 23657 21176 25172 21178
rect 23657 21120 23662 21176
rect 23718 21120 25172 21176
rect 23657 21118 25172 21120
rect 0 21088 800 21118
rect 23657 21115 23723 21118
rect 24372 21088 25172 21118
rect 4469 20704 4785 20705
rect 4469 20640 4475 20704
rect 4539 20640 4555 20704
rect 4619 20640 4635 20704
rect 4699 20640 4715 20704
rect 4779 20640 4785 20704
rect 4469 20639 4785 20640
rect 10196 20704 10512 20705
rect 10196 20640 10202 20704
rect 10266 20640 10282 20704
rect 10346 20640 10362 20704
rect 10426 20640 10442 20704
rect 10506 20640 10512 20704
rect 10196 20639 10512 20640
rect 15923 20704 16239 20705
rect 15923 20640 15929 20704
rect 15993 20640 16009 20704
rect 16073 20640 16089 20704
rect 16153 20640 16169 20704
rect 16233 20640 16239 20704
rect 15923 20639 16239 20640
rect 21650 20704 21966 20705
rect 21650 20640 21656 20704
rect 21720 20640 21736 20704
rect 21800 20640 21816 20704
rect 21880 20640 21896 20704
rect 21960 20640 21966 20704
rect 21650 20639 21966 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 23381 20498 23447 20501
rect 24372 20498 25172 20528
rect 23381 20496 25172 20498
rect 23381 20440 23386 20496
rect 23442 20440 25172 20496
rect 23381 20438 25172 20440
rect 23381 20435 23447 20438
rect 24372 20408 25172 20438
rect 3809 20160 4125 20161
rect 3809 20096 3815 20160
rect 3879 20096 3895 20160
rect 3959 20096 3975 20160
rect 4039 20096 4055 20160
rect 4119 20096 4125 20160
rect 3809 20095 4125 20096
rect 9536 20160 9852 20161
rect 9536 20096 9542 20160
rect 9606 20096 9622 20160
rect 9686 20096 9702 20160
rect 9766 20096 9782 20160
rect 9846 20096 9852 20160
rect 9536 20095 9852 20096
rect 15263 20160 15579 20161
rect 15263 20096 15269 20160
rect 15333 20096 15349 20160
rect 15413 20096 15429 20160
rect 15493 20096 15509 20160
rect 15573 20096 15579 20160
rect 15263 20095 15579 20096
rect 20990 20160 21306 20161
rect 20990 20096 20996 20160
rect 21060 20096 21076 20160
rect 21140 20096 21156 20160
rect 21220 20096 21236 20160
rect 21300 20096 21306 20160
rect 20990 20095 21306 20096
rect 841 19954 907 19957
rect 798 19952 907 19954
rect 798 19896 846 19952
rect 902 19896 907 19952
rect 798 19891 907 19896
rect 798 19848 858 19891
rect 0 19758 858 19848
rect 23657 19818 23723 19821
rect 24372 19818 25172 19848
rect 23657 19816 25172 19818
rect 23657 19760 23662 19816
rect 23718 19760 25172 19816
rect 23657 19758 25172 19760
rect 0 19728 800 19758
rect 23657 19755 23723 19758
rect 24372 19728 25172 19758
rect 4469 19616 4785 19617
rect 4469 19552 4475 19616
rect 4539 19552 4555 19616
rect 4619 19552 4635 19616
rect 4699 19552 4715 19616
rect 4779 19552 4785 19616
rect 4469 19551 4785 19552
rect 10196 19616 10512 19617
rect 10196 19552 10202 19616
rect 10266 19552 10282 19616
rect 10346 19552 10362 19616
rect 10426 19552 10442 19616
rect 10506 19552 10512 19616
rect 10196 19551 10512 19552
rect 15923 19616 16239 19617
rect 15923 19552 15929 19616
rect 15993 19552 16009 19616
rect 16073 19552 16089 19616
rect 16153 19552 16169 19616
rect 16233 19552 16239 19616
rect 15923 19551 16239 19552
rect 21650 19616 21966 19617
rect 21650 19552 21656 19616
rect 21720 19552 21736 19616
rect 21800 19552 21816 19616
rect 21880 19552 21896 19616
rect 21960 19552 21966 19616
rect 21650 19551 21966 19552
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 23381 19138 23447 19141
rect 24372 19138 25172 19168
rect 23381 19136 25172 19138
rect 23381 19080 23386 19136
rect 23442 19080 25172 19136
rect 23381 19078 25172 19080
rect 23381 19075 23447 19078
rect 3809 19072 4125 19073
rect 3809 19008 3815 19072
rect 3879 19008 3895 19072
rect 3959 19008 3975 19072
rect 4039 19008 4055 19072
rect 4119 19008 4125 19072
rect 3809 19007 4125 19008
rect 9536 19072 9852 19073
rect 9536 19008 9542 19072
rect 9606 19008 9622 19072
rect 9686 19008 9702 19072
rect 9766 19008 9782 19072
rect 9846 19008 9852 19072
rect 9536 19007 9852 19008
rect 15263 19072 15579 19073
rect 15263 19008 15269 19072
rect 15333 19008 15349 19072
rect 15413 19008 15429 19072
rect 15493 19008 15509 19072
rect 15573 19008 15579 19072
rect 15263 19007 15579 19008
rect 20990 19072 21306 19073
rect 20990 19008 20996 19072
rect 21060 19008 21076 19072
rect 21140 19008 21156 19072
rect 21220 19008 21236 19072
rect 21300 19008 21306 19072
rect 24372 19048 25172 19078
rect 20990 19007 21306 19008
rect 841 18594 907 18597
rect 798 18592 907 18594
rect 798 18536 846 18592
rect 902 18536 907 18592
rect 798 18531 907 18536
rect 798 18488 858 18531
rect 0 18398 858 18488
rect 4469 18528 4785 18529
rect 4469 18464 4475 18528
rect 4539 18464 4555 18528
rect 4619 18464 4635 18528
rect 4699 18464 4715 18528
rect 4779 18464 4785 18528
rect 4469 18463 4785 18464
rect 10196 18528 10512 18529
rect 10196 18464 10202 18528
rect 10266 18464 10282 18528
rect 10346 18464 10362 18528
rect 10426 18464 10442 18528
rect 10506 18464 10512 18528
rect 10196 18463 10512 18464
rect 15923 18528 16239 18529
rect 15923 18464 15929 18528
rect 15993 18464 16009 18528
rect 16073 18464 16089 18528
rect 16153 18464 16169 18528
rect 16233 18464 16239 18528
rect 15923 18463 16239 18464
rect 21650 18528 21966 18529
rect 21650 18464 21656 18528
rect 21720 18464 21736 18528
rect 21800 18464 21816 18528
rect 21880 18464 21896 18528
rect 21960 18464 21966 18528
rect 21650 18463 21966 18464
rect 23289 18458 23355 18461
rect 24372 18458 25172 18488
rect 23289 18456 25172 18458
rect 23289 18400 23294 18456
rect 23350 18400 25172 18456
rect 23289 18398 25172 18400
rect 0 18368 800 18398
rect 23289 18395 23355 18398
rect 24372 18368 25172 18398
rect 3809 17984 4125 17985
rect 3809 17920 3815 17984
rect 3879 17920 3895 17984
rect 3959 17920 3975 17984
rect 4039 17920 4055 17984
rect 4119 17920 4125 17984
rect 3809 17919 4125 17920
rect 9536 17984 9852 17985
rect 9536 17920 9542 17984
rect 9606 17920 9622 17984
rect 9686 17920 9702 17984
rect 9766 17920 9782 17984
rect 9846 17920 9852 17984
rect 9536 17919 9852 17920
rect 15263 17984 15579 17985
rect 15263 17920 15269 17984
rect 15333 17920 15349 17984
rect 15413 17920 15429 17984
rect 15493 17920 15509 17984
rect 15573 17920 15579 17984
rect 15263 17919 15579 17920
rect 20990 17984 21306 17985
rect 20990 17920 20996 17984
rect 21060 17920 21076 17984
rect 21140 17920 21156 17984
rect 21220 17920 21236 17984
rect 21300 17920 21306 17984
rect 20990 17919 21306 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 23657 17778 23723 17781
rect 24372 17778 25172 17808
rect 23657 17776 25172 17778
rect 23657 17720 23662 17776
rect 23718 17720 25172 17776
rect 23657 17718 25172 17720
rect 23657 17715 23723 17718
rect 24372 17688 25172 17718
rect 4469 17440 4785 17441
rect 4469 17376 4475 17440
rect 4539 17376 4555 17440
rect 4619 17376 4635 17440
rect 4699 17376 4715 17440
rect 4779 17376 4785 17440
rect 4469 17375 4785 17376
rect 10196 17440 10512 17441
rect 10196 17376 10202 17440
rect 10266 17376 10282 17440
rect 10346 17376 10362 17440
rect 10426 17376 10442 17440
rect 10506 17376 10512 17440
rect 10196 17375 10512 17376
rect 15923 17440 16239 17441
rect 15923 17376 15929 17440
rect 15993 17376 16009 17440
rect 16073 17376 16089 17440
rect 16153 17376 16169 17440
rect 16233 17376 16239 17440
rect 15923 17375 16239 17376
rect 21650 17440 21966 17441
rect 21650 17376 21656 17440
rect 21720 17376 21736 17440
rect 21800 17376 21816 17440
rect 21880 17376 21896 17440
rect 21960 17376 21966 17440
rect 21650 17375 21966 17376
rect 841 17234 907 17237
rect 798 17232 907 17234
rect 798 17176 846 17232
rect 902 17176 907 17232
rect 798 17171 907 17176
rect 798 17128 858 17171
rect 0 17038 858 17128
rect 23657 17098 23723 17101
rect 24372 17098 25172 17128
rect 23657 17096 25172 17098
rect 23657 17040 23662 17096
rect 23718 17040 25172 17096
rect 23657 17038 25172 17040
rect 0 17008 800 17038
rect 23657 17035 23723 17038
rect 24372 17008 25172 17038
rect 3809 16896 4125 16897
rect 3809 16832 3815 16896
rect 3879 16832 3895 16896
rect 3959 16832 3975 16896
rect 4039 16832 4055 16896
rect 4119 16832 4125 16896
rect 3809 16831 4125 16832
rect 9536 16896 9852 16897
rect 9536 16832 9542 16896
rect 9606 16832 9622 16896
rect 9686 16832 9702 16896
rect 9766 16832 9782 16896
rect 9846 16832 9852 16896
rect 9536 16831 9852 16832
rect 15263 16896 15579 16897
rect 15263 16832 15269 16896
rect 15333 16832 15349 16896
rect 15413 16832 15429 16896
rect 15493 16832 15509 16896
rect 15573 16832 15579 16896
rect 15263 16831 15579 16832
rect 20990 16896 21306 16897
rect 20990 16832 20996 16896
rect 21060 16832 21076 16896
rect 21140 16832 21156 16896
rect 21220 16832 21236 16896
rect 21300 16832 21306 16896
rect 20990 16831 21306 16832
rect 841 16554 907 16557
rect 798 16552 907 16554
rect 798 16496 846 16552
rect 902 16496 907 16552
rect 798 16491 907 16496
rect 22001 16554 22067 16557
rect 23197 16554 23263 16557
rect 22001 16552 23263 16554
rect 22001 16496 22006 16552
rect 22062 16496 23202 16552
rect 23258 16496 23263 16552
rect 22001 16494 23263 16496
rect 22001 16491 22067 16494
rect 23197 16491 23263 16494
rect 798 16448 858 16491
rect 0 16358 858 16448
rect 23657 16418 23723 16421
rect 24372 16418 25172 16448
rect 23657 16416 25172 16418
rect 23657 16360 23662 16416
rect 23718 16360 25172 16416
rect 23657 16358 25172 16360
rect 0 16328 800 16358
rect 23657 16355 23723 16358
rect 4469 16352 4785 16353
rect 4469 16288 4475 16352
rect 4539 16288 4555 16352
rect 4619 16288 4635 16352
rect 4699 16288 4715 16352
rect 4779 16288 4785 16352
rect 4469 16287 4785 16288
rect 10196 16352 10512 16353
rect 10196 16288 10202 16352
rect 10266 16288 10282 16352
rect 10346 16288 10362 16352
rect 10426 16288 10442 16352
rect 10506 16288 10512 16352
rect 10196 16287 10512 16288
rect 15923 16352 16239 16353
rect 15923 16288 15929 16352
rect 15993 16288 16009 16352
rect 16073 16288 16089 16352
rect 16153 16288 16169 16352
rect 16233 16288 16239 16352
rect 15923 16287 16239 16288
rect 21650 16352 21966 16353
rect 21650 16288 21656 16352
rect 21720 16288 21736 16352
rect 21800 16288 21816 16352
rect 21880 16288 21896 16352
rect 21960 16288 21966 16352
rect 24372 16328 25172 16358
rect 21650 16287 21966 16288
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 3809 15808 4125 15809
rect 3809 15744 3815 15808
rect 3879 15744 3895 15808
rect 3959 15744 3975 15808
rect 4039 15744 4055 15808
rect 4119 15744 4125 15808
rect 3809 15743 4125 15744
rect 9536 15808 9852 15809
rect 9536 15744 9542 15808
rect 9606 15744 9622 15808
rect 9686 15744 9702 15808
rect 9766 15744 9782 15808
rect 9846 15744 9852 15808
rect 9536 15743 9852 15744
rect 15263 15808 15579 15809
rect 15263 15744 15269 15808
rect 15333 15744 15349 15808
rect 15413 15744 15429 15808
rect 15493 15744 15509 15808
rect 15573 15744 15579 15808
rect 15263 15743 15579 15744
rect 20990 15808 21306 15809
rect 20990 15744 20996 15808
rect 21060 15744 21076 15808
rect 21140 15744 21156 15808
rect 21220 15744 21236 15808
rect 21300 15744 21306 15808
rect 20990 15743 21306 15744
rect 23657 15738 23723 15741
rect 24372 15738 25172 15768
rect 23657 15736 25172 15738
rect 23657 15680 23662 15736
rect 23718 15680 25172 15736
rect 23657 15678 25172 15680
rect 0 15648 800 15678
rect 23657 15675 23723 15678
rect 24372 15648 25172 15678
rect 4469 15264 4785 15265
rect 4469 15200 4475 15264
rect 4539 15200 4555 15264
rect 4619 15200 4635 15264
rect 4699 15200 4715 15264
rect 4779 15200 4785 15264
rect 4469 15199 4785 15200
rect 10196 15264 10512 15265
rect 10196 15200 10202 15264
rect 10266 15200 10282 15264
rect 10346 15200 10362 15264
rect 10426 15200 10442 15264
rect 10506 15200 10512 15264
rect 10196 15199 10512 15200
rect 15923 15264 16239 15265
rect 15923 15200 15929 15264
rect 15993 15200 16009 15264
rect 16073 15200 16089 15264
rect 16153 15200 16169 15264
rect 16233 15200 16239 15264
rect 15923 15199 16239 15200
rect 21650 15264 21966 15265
rect 21650 15200 21656 15264
rect 21720 15200 21736 15264
rect 21800 15200 21816 15264
rect 21880 15200 21896 15264
rect 21960 15200 21966 15264
rect 21650 15199 21966 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 23381 15058 23447 15061
rect 24372 15058 25172 15088
rect 23381 15056 25172 15058
rect 23381 15000 23386 15056
rect 23442 15000 25172 15056
rect 23381 14998 25172 15000
rect 23381 14995 23447 14998
rect 24372 14968 25172 14998
rect 3809 14720 4125 14721
rect 3809 14656 3815 14720
rect 3879 14656 3895 14720
rect 3959 14656 3975 14720
rect 4039 14656 4055 14720
rect 4119 14656 4125 14720
rect 3809 14655 4125 14656
rect 9536 14720 9852 14721
rect 9536 14656 9542 14720
rect 9606 14656 9622 14720
rect 9686 14656 9702 14720
rect 9766 14656 9782 14720
rect 9846 14656 9852 14720
rect 9536 14655 9852 14656
rect 15263 14720 15579 14721
rect 15263 14656 15269 14720
rect 15333 14656 15349 14720
rect 15413 14656 15429 14720
rect 15493 14656 15509 14720
rect 15573 14656 15579 14720
rect 15263 14655 15579 14656
rect 20990 14720 21306 14721
rect 20990 14656 20996 14720
rect 21060 14656 21076 14720
rect 21140 14656 21156 14720
rect 21220 14656 21236 14720
rect 21300 14656 21306 14720
rect 20990 14655 21306 14656
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 23657 14378 23723 14381
rect 24372 14378 25172 14408
rect 23657 14376 25172 14378
rect 23657 14320 23662 14376
rect 23718 14320 25172 14376
rect 23657 14318 25172 14320
rect 0 14288 800 14318
rect 23657 14315 23723 14318
rect 24372 14288 25172 14318
rect 4469 14176 4785 14177
rect 4469 14112 4475 14176
rect 4539 14112 4555 14176
rect 4619 14112 4635 14176
rect 4699 14112 4715 14176
rect 4779 14112 4785 14176
rect 4469 14111 4785 14112
rect 10196 14176 10512 14177
rect 10196 14112 10202 14176
rect 10266 14112 10282 14176
rect 10346 14112 10362 14176
rect 10426 14112 10442 14176
rect 10506 14112 10512 14176
rect 10196 14111 10512 14112
rect 15923 14176 16239 14177
rect 15923 14112 15929 14176
rect 15993 14112 16009 14176
rect 16073 14112 16089 14176
rect 16153 14112 16169 14176
rect 16233 14112 16239 14176
rect 15923 14111 16239 14112
rect 21650 14176 21966 14177
rect 21650 14112 21656 14176
rect 21720 14112 21736 14176
rect 21800 14112 21816 14176
rect 21880 14112 21896 14176
rect 21960 14112 21966 14176
rect 21650 14111 21966 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 23381 13698 23447 13701
rect 24372 13698 25172 13728
rect 23381 13696 25172 13698
rect 23381 13640 23386 13696
rect 23442 13640 25172 13696
rect 23381 13638 25172 13640
rect 23381 13635 23447 13638
rect 3809 13632 4125 13633
rect 3809 13568 3815 13632
rect 3879 13568 3895 13632
rect 3959 13568 3975 13632
rect 4039 13568 4055 13632
rect 4119 13568 4125 13632
rect 3809 13567 4125 13568
rect 9536 13632 9852 13633
rect 9536 13568 9542 13632
rect 9606 13568 9622 13632
rect 9686 13568 9702 13632
rect 9766 13568 9782 13632
rect 9846 13568 9852 13632
rect 9536 13567 9852 13568
rect 15263 13632 15579 13633
rect 15263 13568 15269 13632
rect 15333 13568 15349 13632
rect 15413 13568 15429 13632
rect 15493 13568 15509 13632
rect 15573 13568 15579 13632
rect 15263 13567 15579 13568
rect 20990 13632 21306 13633
rect 20990 13568 20996 13632
rect 21060 13568 21076 13632
rect 21140 13568 21156 13632
rect 21220 13568 21236 13632
rect 21300 13568 21306 13632
rect 24372 13608 25172 13638
rect 20990 13567 21306 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 4469 13088 4785 13089
rect 4469 13024 4475 13088
rect 4539 13024 4555 13088
rect 4619 13024 4635 13088
rect 4699 13024 4715 13088
rect 4779 13024 4785 13088
rect 4469 13023 4785 13024
rect 10196 13088 10512 13089
rect 10196 13024 10202 13088
rect 10266 13024 10282 13088
rect 10346 13024 10362 13088
rect 10426 13024 10442 13088
rect 10506 13024 10512 13088
rect 10196 13023 10512 13024
rect 15923 13088 16239 13089
rect 15923 13024 15929 13088
rect 15993 13024 16009 13088
rect 16073 13024 16089 13088
rect 16153 13024 16169 13088
rect 16233 13024 16239 13088
rect 15923 13023 16239 13024
rect 21650 13088 21966 13089
rect 21650 13024 21656 13088
rect 21720 13024 21736 13088
rect 21800 13024 21816 13088
rect 21880 13024 21896 13088
rect 21960 13024 21966 13088
rect 21650 13023 21966 13024
rect 23657 13018 23723 13021
rect 24372 13018 25172 13048
rect 23657 13016 25172 13018
rect 23657 12960 23662 13016
rect 23718 12960 25172 13016
rect 23657 12958 25172 12960
rect 0 12928 800 12958
rect 23657 12955 23723 12958
rect 24372 12928 25172 12958
rect 3809 12544 4125 12545
rect 3809 12480 3815 12544
rect 3879 12480 3895 12544
rect 3959 12480 3975 12544
rect 4039 12480 4055 12544
rect 4119 12480 4125 12544
rect 3809 12479 4125 12480
rect 9536 12544 9852 12545
rect 9536 12480 9542 12544
rect 9606 12480 9622 12544
rect 9686 12480 9702 12544
rect 9766 12480 9782 12544
rect 9846 12480 9852 12544
rect 9536 12479 9852 12480
rect 15263 12544 15579 12545
rect 15263 12480 15269 12544
rect 15333 12480 15349 12544
rect 15413 12480 15429 12544
rect 15493 12480 15509 12544
rect 15573 12480 15579 12544
rect 15263 12479 15579 12480
rect 20990 12544 21306 12545
rect 20990 12480 20996 12544
rect 21060 12480 21076 12544
rect 21140 12480 21156 12544
rect 21220 12480 21236 12544
rect 21300 12480 21306 12544
rect 20990 12479 21306 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 23381 12338 23447 12341
rect 24372 12338 25172 12368
rect 23381 12336 25172 12338
rect 23381 12280 23386 12336
rect 23442 12280 25172 12336
rect 23381 12278 25172 12280
rect 23381 12275 23447 12278
rect 24372 12248 25172 12278
rect 4469 12000 4785 12001
rect 4469 11936 4475 12000
rect 4539 11936 4555 12000
rect 4619 11936 4635 12000
rect 4699 11936 4715 12000
rect 4779 11936 4785 12000
rect 4469 11935 4785 11936
rect 10196 12000 10512 12001
rect 10196 11936 10202 12000
rect 10266 11936 10282 12000
rect 10346 11936 10362 12000
rect 10426 11936 10442 12000
rect 10506 11936 10512 12000
rect 10196 11935 10512 11936
rect 15923 12000 16239 12001
rect 15923 11936 15929 12000
rect 15993 11936 16009 12000
rect 16073 11936 16089 12000
rect 16153 11936 16169 12000
rect 16233 11936 16239 12000
rect 15923 11935 16239 11936
rect 21650 12000 21966 12001
rect 21650 11936 21656 12000
rect 21720 11936 21736 12000
rect 21800 11936 21816 12000
rect 21880 11936 21896 12000
rect 21960 11936 21966 12000
rect 21650 11935 21966 11936
rect 841 11794 907 11797
rect 798 11792 907 11794
rect 798 11736 846 11792
rect 902 11736 907 11792
rect 798 11731 907 11736
rect 798 11688 858 11731
rect 0 11598 858 11688
rect 23657 11658 23723 11661
rect 24372 11658 25172 11688
rect 23657 11656 25172 11658
rect 23657 11600 23662 11656
rect 23718 11600 25172 11656
rect 23657 11598 25172 11600
rect 0 11568 800 11598
rect 23657 11595 23723 11598
rect 24372 11568 25172 11598
rect 3809 11456 4125 11457
rect 3809 11392 3815 11456
rect 3879 11392 3895 11456
rect 3959 11392 3975 11456
rect 4039 11392 4055 11456
rect 4119 11392 4125 11456
rect 3809 11391 4125 11392
rect 9536 11456 9852 11457
rect 9536 11392 9542 11456
rect 9606 11392 9622 11456
rect 9686 11392 9702 11456
rect 9766 11392 9782 11456
rect 9846 11392 9852 11456
rect 9536 11391 9852 11392
rect 15263 11456 15579 11457
rect 15263 11392 15269 11456
rect 15333 11392 15349 11456
rect 15413 11392 15429 11456
rect 15493 11392 15509 11456
rect 15573 11392 15579 11456
rect 15263 11391 15579 11392
rect 20990 11456 21306 11457
rect 20990 11392 20996 11456
rect 21060 11392 21076 11456
rect 21140 11392 21156 11456
rect 21220 11392 21236 11456
rect 21300 11392 21306 11456
rect 20990 11391 21306 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 23381 10978 23447 10981
rect 24372 10978 25172 11008
rect 23381 10976 25172 10978
rect 23381 10920 23386 10976
rect 23442 10920 25172 10976
rect 23381 10918 25172 10920
rect 23381 10915 23447 10918
rect 4469 10912 4785 10913
rect 4469 10848 4475 10912
rect 4539 10848 4555 10912
rect 4619 10848 4635 10912
rect 4699 10848 4715 10912
rect 4779 10848 4785 10912
rect 4469 10847 4785 10848
rect 10196 10912 10512 10913
rect 10196 10848 10202 10912
rect 10266 10848 10282 10912
rect 10346 10848 10362 10912
rect 10426 10848 10442 10912
rect 10506 10848 10512 10912
rect 10196 10847 10512 10848
rect 15923 10912 16239 10913
rect 15923 10848 15929 10912
rect 15993 10848 16009 10912
rect 16073 10848 16089 10912
rect 16153 10848 16169 10912
rect 16233 10848 16239 10912
rect 15923 10847 16239 10848
rect 21650 10912 21966 10913
rect 21650 10848 21656 10912
rect 21720 10848 21736 10912
rect 21800 10848 21816 10912
rect 21880 10848 21896 10912
rect 21960 10848 21966 10912
rect 24372 10888 25172 10918
rect 21650 10847 21966 10848
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 3809 10368 4125 10369
rect 3809 10304 3815 10368
rect 3879 10304 3895 10368
rect 3959 10304 3975 10368
rect 4039 10304 4055 10368
rect 4119 10304 4125 10368
rect 3809 10303 4125 10304
rect 9536 10368 9852 10369
rect 9536 10304 9542 10368
rect 9606 10304 9622 10368
rect 9686 10304 9702 10368
rect 9766 10304 9782 10368
rect 9846 10304 9852 10368
rect 9536 10303 9852 10304
rect 15263 10368 15579 10369
rect 15263 10304 15269 10368
rect 15333 10304 15349 10368
rect 15413 10304 15429 10368
rect 15493 10304 15509 10368
rect 15573 10304 15579 10368
rect 15263 10303 15579 10304
rect 20990 10368 21306 10369
rect 20990 10304 20996 10368
rect 21060 10304 21076 10368
rect 21140 10304 21156 10368
rect 21220 10304 21236 10368
rect 21300 10304 21306 10368
rect 20990 10303 21306 10304
rect 23657 10298 23723 10301
rect 24372 10298 25172 10328
rect 23657 10296 25172 10298
rect 23657 10240 23662 10296
rect 23718 10240 25172 10296
rect 23657 10238 25172 10240
rect 0 10208 800 10238
rect 23657 10235 23723 10238
rect 24372 10208 25172 10238
rect 4469 9824 4785 9825
rect 4469 9760 4475 9824
rect 4539 9760 4555 9824
rect 4619 9760 4635 9824
rect 4699 9760 4715 9824
rect 4779 9760 4785 9824
rect 4469 9759 4785 9760
rect 10196 9824 10512 9825
rect 10196 9760 10202 9824
rect 10266 9760 10282 9824
rect 10346 9760 10362 9824
rect 10426 9760 10442 9824
rect 10506 9760 10512 9824
rect 10196 9759 10512 9760
rect 15923 9824 16239 9825
rect 15923 9760 15929 9824
rect 15993 9760 16009 9824
rect 16073 9760 16089 9824
rect 16153 9760 16169 9824
rect 16233 9760 16239 9824
rect 15923 9759 16239 9760
rect 21650 9824 21966 9825
rect 21650 9760 21656 9824
rect 21720 9760 21736 9824
rect 21800 9760 21816 9824
rect 21880 9760 21896 9824
rect 21960 9760 21966 9824
rect 21650 9759 21966 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 23657 9618 23723 9621
rect 24372 9618 25172 9648
rect 23657 9616 25172 9618
rect 23657 9560 23662 9616
rect 23718 9560 25172 9616
rect 23657 9558 25172 9560
rect 23657 9555 23723 9558
rect 24372 9528 25172 9558
rect 3809 9280 4125 9281
rect 3809 9216 3815 9280
rect 3879 9216 3895 9280
rect 3959 9216 3975 9280
rect 4039 9216 4055 9280
rect 4119 9216 4125 9280
rect 3809 9215 4125 9216
rect 9536 9280 9852 9281
rect 9536 9216 9542 9280
rect 9606 9216 9622 9280
rect 9686 9216 9702 9280
rect 9766 9216 9782 9280
rect 9846 9216 9852 9280
rect 9536 9215 9852 9216
rect 15263 9280 15579 9281
rect 15263 9216 15269 9280
rect 15333 9216 15349 9280
rect 15413 9216 15429 9280
rect 15493 9216 15509 9280
rect 15573 9216 15579 9280
rect 15263 9215 15579 9216
rect 20990 9280 21306 9281
rect 20990 9216 20996 9280
rect 21060 9216 21076 9280
rect 21140 9216 21156 9280
rect 21220 9216 21236 9280
rect 21300 9216 21306 9280
rect 20990 9215 21306 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 23657 8938 23723 8941
rect 24372 8938 25172 8968
rect 23657 8936 25172 8938
rect 23657 8880 23662 8936
rect 23718 8880 25172 8936
rect 23657 8878 25172 8880
rect 0 8848 800 8878
rect 23657 8875 23723 8878
rect 24372 8848 25172 8878
rect 4469 8736 4785 8737
rect 4469 8672 4475 8736
rect 4539 8672 4555 8736
rect 4619 8672 4635 8736
rect 4699 8672 4715 8736
rect 4779 8672 4785 8736
rect 4469 8671 4785 8672
rect 10196 8736 10512 8737
rect 10196 8672 10202 8736
rect 10266 8672 10282 8736
rect 10346 8672 10362 8736
rect 10426 8672 10442 8736
rect 10506 8672 10512 8736
rect 10196 8671 10512 8672
rect 15923 8736 16239 8737
rect 15923 8672 15929 8736
rect 15993 8672 16009 8736
rect 16073 8672 16089 8736
rect 16153 8672 16169 8736
rect 16233 8672 16239 8736
rect 15923 8671 16239 8672
rect 21650 8736 21966 8737
rect 21650 8672 21656 8736
rect 21720 8672 21736 8736
rect 21800 8672 21816 8736
rect 21880 8672 21896 8736
rect 21960 8672 21966 8736
rect 21650 8671 21966 8672
rect 23381 8258 23447 8261
rect 24372 8258 25172 8288
rect 23381 8256 25172 8258
rect 23381 8200 23386 8256
rect 23442 8200 25172 8256
rect 23381 8198 25172 8200
rect 23381 8195 23447 8198
rect 3809 8192 4125 8193
rect 3809 8128 3815 8192
rect 3879 8128 3895 8192
rect 3959 8128 3975 8192
rect 4039 8128 4055 8192
rect 4119 8128 4125 8192
rect 3809 8127 4125 8128
rect 9536 8192 9852 8193
rect 9536 8128 9542 8192
rect 9606 8128 9622 8192
rect 9686 8128 9702 8192
rect 9766 8128 9782 8192
rect 9846 8128 9852 8192
rect 9536 8127 9852 8128
rect 15263 8192 15579 8193
rect 15263 8128 15269 8192
rect 15333 8128 15349 8192
rect 15413 8128 15429 8192
rect 15493 8128 15509 8192
rect 15573 8128 15579 8192
rect 15263 8127 15579 8128
rect 20990 8192 21306 8193
rect 20990 8128 20996 8192
rect 21060 8128 21076 8192
rect 21140 8128 21156 8192
rect 21220 8128 21236 8192
rect 21300 8128 21306 8192
rect 24372 8168 25172 8198
rect 20990 8127 21306 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4469 7648 4785 7649
rect 4469 7584 4475 7648
rect 4539 7584 4555 7648
rect 4619 7584 4635 7648
rect 4699 7584 4715 7648
rect 4779 7584 4785 7648
rect 4469 7583 4785 7584
rect 10196 7648 10512 7649
rect 10196 7584 10202 7648
rect 10266 7584 10282 7648
rect 10346 7584 10362 7648
rect 10426 7584 10442 7648
rect 10506 7584 10512 7648
rect 10196 7583 10512 7584
rect 15923 7648 16239 7649
rect 15923 7584 15929 7648
rect 15993 7584 16009 7648
rect 16073 7584 16089 7648
rect 16153 7584 16169 7648
rect 16233 7584 16239 7648
rect 15923 7583 16239 7584
rect 21650 7648 21966 7649
rect 21650 7584 21656 7648
rect 21720 7584 21736 7648
rect 21800 7584 21816 7648
rect 21880 7584 21896 7648
rect 21960 7584 21966 7648
rect 21650 7583 21966 7584
rect 23657 7578 23723 7581
rect 24372 7578 25172 7608
rect 23657 7576 25172 7578
rect 23657 7520 23662 7576
rect 23718 7520 25172 7576
rect 23657 7518 25172 7520
rect 0 7488 800 7518
rect 23657 7515 23723 7518
rect 24372 7488 25172 7518
rect 3809 7104 4125 7105
rect 3809 7040 3815 7104
rect 3879 7040 3895 7104
rect 3959 7040 3975 7104
rect 4039 7040 4055 7104
rect 4119 7040 4125 7104
rect 3809 7039 4125 7040
rect 9536 7104 9852 7105
rect 9536 7040 9542 7104
rect 9606 7040 9622 7104
rect 9686 7040 9702 7104
rect 9766 7040 9782 7104
rect 9846 7040 9852 7104
rect 9536 7039 9852 7040
rect 15263 7104 15579 7105
rect 15263 7040 15269 7104
rect 15333 7040 15349 7104
rect 15413 7040 15429 7104
rect 15493 7040 15509 7104
rect 15573 7040 15579 7104
rect 15263 7039 15579 7040
rect 20990 7104 21306 7105
rect 20990 7040 20996 7104
rect 21060 7040 21076 7104
rect 21140 7040 21156 7104
rect 21220 7040 21236 7104
rect 21300 7040 21306 7104
rect 20990 7039 21306 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 23657 6898 23723 6901
rect 24372 6898 25172 6928
rect 23657 6896 25172 6898
rect 23657 6840 23662 6896
rect 23718 6840 25172 6896
rect 23657 6838 25172 6840
rect 23657 6835 23723 6838
rect 24372 6808 25172 6838
rect 4469 6560 4785 6561
rect 4469 6496 4475 6560
rect 4539 6496 4555 6560
rect 4619 6496 4635 6560
rect 4699 6496 4715 6560
rect 4779 6496 4785 6560
rect 4469 6495 4785 6496
rect 10196 6560 10512 6561
rect 10196 6496 10202 6560
rect 10266 6496 10282 6560
rect 10346 6496 10362 6560
rect 10426 6496 10442 6560
rect 10506 6496 10512 6560
rect 10196 6495 10512 6496
rect 15923 6560 16239 6561
rect 15923 6496 15929 6560
rect 15993 6496 16009 6560
rect 16073 6496 16089 6560
rect 16153 6496 16169 6560
rect 16233 6496 16239 6560
rect 15923 6495 16239 6496
rect 21650 6560 21966 6561
rect 21650 6496 21656 6560
rect 21720 6496 21736 6560
rect 21800 6496 21816 6560
rect 21880 6496 21896 6560
rect 21960 6496 21966 6560
rect 21650 6495 21966 6496
rect 23657 6218 23723 6221
rect 24372 6218 25172 6248
rect 23657 6216 25172 6218
rect 23657 6160 23662 6216
rect 23718 6160 25172 6216
rect 23657 6158 25172 6160
rect 23657 6155 23723 6158
rect 24372 6128 25172 6158
rect 3809 6016 4125 6017
rect 3809 5952 3815 6016
rect 3879 5952 3895 6016
rect 3959 5952 3975 6016
rect 4039 5952 4055 6016
rect 4119 5952 4125 6016
rect 3809 5951 4125 5952
rect 9536 6016 9852 6017
rect 9536 5952 9542 6016
rect 9606 5952 9622 6016
rect 9686 5952 9702 6016
rect 9766 5952 9782 6016
rect 9846 5952 9852 6016
rect 9536 5951 9852 5952
rect 15263 6016 15579 6017
rect 15263 5952 15269 6016
rect 15333 5952 15349 6016
rect 15413 5952 15429 6016
rect 15493 5952 15509 6016
rect 15573 5952 15579 6016
rect 15263 5951 15579 5952
rect 20990 6016 21306 6017
rect 20990 5952 20996 6016
rect 21060 5952 21076 6016
rect 21140 5952 21156 6016
rect 21220 5952 21236 6016
rect 21300 5952 21306 6016
rect 20990 5951 21306 5952
rect 23381 5538 23447 5541
rect 24372 5538 25172 5568
rect 23381 5536 25172 5538
rect 23381 5480 23386 5536
rect 23442 5480 25172 5536
rect 23381 5478 25172 5480
rect 23381 5475 23447 5478
rect 4469 5472 4785 5473
rect 4469 5408 4475 5472
rect 4539 5408 4555 5472
rect 4619 5408 4635 5472
rect 4699 5408 4715 5472
rect 4779 5408 4785 5472
rect 4469 5407 4785 5408
rect 10196 5472 10512 5473
rect 10196 5408 10202 5472
rect 10266 5408 10282 5472
rect 10346 5408 10362 5472
rect 10426 5408 10442 5472
rect 10506 5408 10512 5472
rect 10196 5407 10512 5408
rect 15923 5472 16239 5473
rect 15923 5408 15929 5472
rect 15993 5408 16009 5472
rect 16073 5408 16089 5472
rect 16153 5408 16169 5472
rect 16233 5408 16239 5472
rect 15923 5407 16239 5408
rect 21650 5472 21966 5473
rect 21650 5408 21656 5472
rect 21720 5408 21736 5472
rect 21800 5408 21816 5472
rect 21880 5408 21896 5472
rect 21960 5408 21966 5472
rect 24372 5448 25172 5478
rect 21650 5407 21966 5408
rect 3809 4928 4125 4929
rect 3809 4864 3815 4928
rect 3879 4864 3895 4928
rect 3959 4864 3975 4928
rect 4039 4864 4055 4928
rect 4119 4864 4125 4928
rect 3809 4863 4125 4864
rect 9536 4928 9852 4929
rect 9536 4864 9542 4928
rect 9606 4864 9622 4928
rect 9686 4864 9702 4928
rect 9766 4864 9782 4928
rect 9846 4864 9852 4928
rect 9536 4863 9852 4864
rect 15263 4928 15579 4929
rect 15263 4864 15269 4928
rect 15333 4864 15349 4928
rect 15413 4864 15429 4928
rect 15493 4864 15509 4928
rect 15573 4864 15579 4928
rect 15263 4863 15579 4864
rect 20990 4928 21306 4929
rect 20990 4864 20996 4928
rect 21060 4864 21076 4928
rect 21140 4864 21156 4928
rect 21220 4864 21236 4928
rect 21300 4864 21306 4928
rect 20990 4863 21306 4864
rect 23657 4858 23723 4861
rect 24372 4858 25172 4888
rect 23657 4856 25172 4858
rect 23657 4800 23662 4856
rect 23718 4800 25172 4856
rect 23657 4798 25172 4800
rect 23657 4795 23723 4798
rect 24372 4768 25172 4798
rect 4469 4384 4785 4385
rect 4469 4320 4475 4384
rect 4539 4320 4555 4384
rect 4619 4320 4635 4384
rect 4699 4320 4715 4384
rect 4779 4320 4785 4384
rect 4469 4319 4785 4320
rect 10196 4384 10512 4385
rect 10196 4320 10202 4384
rect 10266 4320 10282 4384
rect 10346 4320 10362 4384
rect 10426 4320 10442 4384
rect 10506 4320 10512 4384
rect 10196 4319 10512 4320
rect 15923 4384 16239 4385
rect 15923 4320 15929 4384
rect 15993 4320 16009 4384
rect 16073 4320 16089 4384
rect 16153 4320 16169 4384
rect 16233 4320 16239 4384
rect 15923 4319 16239 4320
rect 21650 4384 21966 4385
rect 21650 4320 21656 4384
rect 21720 4320 21736 4384
rect 21800 4320 21816 4384
rect 21880 4320 21896 4384
rect 21960 4320 21966 4384
rect 21650 4319 21966 4320
rect 23657 4178 23723 4181
rect 24372 4178 25172 4208
rect 23657 4176 25172 4178
rect 23657 4120 23662 4176
rect 23718 4120 25172 4176
rect 23657 4118 25172 4120
rect 23657 4115 23723 4118
rect 24372 4088 25172 4118
rect 3809 3840 4125 3841
rect 3809 3776 3815 3840
rect 3879 3776 3895 3840
rect 3959 3776 3975 3840
rect 4039 3776 4055 3840
rect 4119 3776 4125 3840
rect 3809 3775 4125 3776
rect 9536 3840 9852 3841
rect 9536 3776 9542 3840
rect 9606 3776 9622 3840
rect 9686 3776 9702 3840
rect 9766 3776 9782 3840
rect 9846 3776 9852 3840
rect 9536 3775 9852 3776
rect 15263 3840 15579 3841
rect 15263 3776 15269 3840
rect 15333 3776 15349 3840
rect 15413 3776 15429 3840
rect 15493 3776 15509 3840
rect 15573 3776 15579 3840
rect 15263 3775 15579 3776
rect 20990 3840 21306 3841
rect 20990 3776 20996 3840
rect 21060 3776 21076 3840
rect 21140 3776 21156 3840
rect 21220 3776 21236 3840
rect 21300 3776 21306 3840
rect 20990 3775 21306 3776
rect 23657 3498 23723 3501
rect 24372 3498 25172 3528
rect 23657 3496 25172 3498
rect 23657 3440 23662 3496
rect 23718 3440 25172 3496
rect 23657 3438 25172 3440
rect 23657 3435 23723 3438
rect 24372 3408 25172 3438
rect 4469 3296 4785 3297
rect 4469 3232 4475 3296
rect 4539 3232 4555 3296
rect 4619 3232 4635 3296
rect 4699 3232 4715 3296
rect 4779 3232 4785 3296
rect 4469 3231 4785 3232
rect 10196 3296 10512 3297
rect 10196 3232 10202 3296
rect 10266 3232 10282 3296
rect 10346 3232 10362 3296
rect 10426 3232 10442 3296
rect 10506 3232 10512 3296
rect 10196 3231 10512 3232
rect 15923 3296 16239 3297
rect 15923 3232 15929 3296
rect 15993 3232 16009 3296
rect 16073 3232 16089 3296
rect 16153 3232 16169 3296
rect 16233 3232 16239 3296
rect 15923 3231 16239 3232
rect 21650 3296 21966 3297
rect 21650 3232 21656 3296
rect 21720 3232 21736 3296
rect 21800 3232 21816 3296
rect 21880 3232 21896 3296
rect 21960 3232 21966 3296
rect 21650 3231 21966 3232
rect 23657 2818 23723 2821
rect 24372 2818 25172 2848
rect 23657 2816 25172 2818
rect 23657 2760 23662 2816
rect 23718 2760 25172 2816
rect 23657 2758 25172 2760
rect 23657 2755 23723 2758
rect 3809 2752 4125 2753
rect 3809 2688 3815 2752
rect 3879 2688 3895 2752
rect 3959 2688 3975 2752
rect 4039 2688 4055 2752
rect 4119 2688 4125 2752
rect 3809 2687 4125 2688
rect 9536 2752 9852 2753
rect 9536 2688 9542 2752
rect 9606 2688 9622 2752
rect 9686 2688 9702 2752
rect 9766 2688 9782 2752
rect 9846 2688 9852 2752
rect 9536 2687 9852 2688
rect 15263 2752 15579 2753
rect 15263 2688 15269 2752
rect 15333 2688 15349 2752
rect 15413 2688 15429 2752
rect 15493 2688 15509 2752
rect 15573 2688 15579 2752
rect 15263 2687 15579 2688
rect 20990 2752 21306 2753
rect 20990 2688 20996 2752
rect 21060 2688 21076 2752
rect 21140 2688 21156 2752
rect 21220 2688 21236 2752
rect 21300 2688 21306 2752
rect 24372 2728 25172 2758
rect 20990 2687 21306 2688
rect 4469 2208 4785 2209
rect 4469 2144 4475 2208
rect 4539 2144 4555 2208
rect 4619 2144 4635 2208
rect 4699 2144 4715 2208
rect 4779 2144 4785 2208
rect 4469 2143 4785 2144
rect 10196 2208 10512 2209
rect 10196 2144 10202 2208
rect 10266 2144 10282 2208
rect 10346 2144 10362 2208
rect 10426 2144 10442 2208
rect 10506 2144 10512 2208
rect 10196 2143 10512 2144
rect 15923 2208 16239 2209
rect 15923 2144 15929 2208
rect 15993 2144 16009 2208
rect 16073 2144 16089 2208
rect 16153 2144 16169 2208
rect 16233 2144 16239 2208
rect 15923 2143 16239 2144
rect 21650 2208 21966 2209
rect 21650 2144 21656 2208
rect 21720 2144 21736 2208
rect 21800 2144 21816 2208
rect 21880 2144 21896 2208
rect 21960 2144 21966 2208
rect 21650 2143 21966 2144
<< via3 >>
rect 4475 25052 4539 25056
rect 4475 24996 4479 25052
rect 4479 24996 4535 25052
rect 4535 24996 4539 25052
rect 4475 24992 4539 24996
rect 4555 25052 4619 25056
rect 4555 24996 4559 25052
rect 4559 24996 4615 25052
rect 4615 24996 4619 25052
rect 4555 24992 4619 24996
rect 4635 25052 4699 25056
rect 4635 24996 4639 25052
rect 4639 24996 4695 25052
rect 4695 24996 4699 25052
rect 4635 24992 4699 24996
rect 4715 25052 4779 25056
rect 4715 24996 4719 25052
rect 4719 24996 4775 25052
rect 4775 24996 4779 25052
rect 4715 24992 4779 24996
rect 10202 25052 10266 25056
rect 10202 24996 10206 25052
rect 10206 24996 10262 25052
rect 10262 24996 10266 25052
rect 10202 24992 10266 24996
rect 10282 25052 10346 25056
rect 10282 24996 10286 25052
rect 10286 24996 10342 25052
rect 10342 24996 10346 25052
rect 10282 24992 10346 24996
rect 10362 25052 10426 25056
rect 10362 24996 10366 25052
rect 10366 24996 10422 25052
rect 10422 24996 10426 25052
rect 10362 24992 10426 24996
rect 10442 25052 10506 25056
rect 10442 24996 10446 25052
rect 10446 24996 10502 25052
rect 10502 24996 10506 25052
rect 10442 24992 10506 24996
rect 15929 25052 15993 25056
rect 15929 24996 15933 25052
rect 15933 24996 15989 25052
rect 15989 24996 15993 25052
rect 15929 24992 15993 24996
rect 16009 25052 16073 25056
rect 16009 24996 16013 25052
rect 16013 24996 16069 25052
rect 16069 24996 16073 25052
rect 16009 24992 16073 24996
rect 16089 25052 16153 25056
rect 16089 24996 16093 25052
rect 16093 24996 16149 25052
rect 16149 24996 16153 25052
rect 16089 24992 16153 24996
rect 16169 25052 16233 25056
rect 16169 24996 16173 25052
rect 16173 24996 16229 25052
rect 16229 24996 16233 25052
rect 16169 24992 16233 24996
rect 21656 25052 21720 25056
rect 21656 24996 21660 25052
rect 21660 24996 21716 25052
rect 21716 24996 21720 25052
rect 21656 24992 21720 24996
rect 21736 25052 21800 25056
rect 21736 24996 21740 25052
rect 21740 24996 21796 25052
rect 21796 24996 21800 25052
rect 21736 24992 21800 24996
rect 21816 25052 21880 25056
rect 21816 24996 21820 25052
rect 21820 24996 21876 25052
rect 21876 24996 21880 25052
rect 21816 24992 21880 24996
rect 21896 25052 21960 25056
rect 21896 24996 21900 25052
rect 21900 24996 21956 25052
rect 21956 24996 21960 25052
rect 21896 24992 21960 24996
rect 3815 24508 3879 24512
rect 3815 24452 3819 24508
rect 3819 24452 3875 24508
rect 3875 24452 3879 24508
rect 3815 24448 3879 24452
rect 3895 24508 3959 24512
rect 3895 24452 3899 24508
rect 3899 24452 3955 24508
rect 3955 24452 3959 24508
rect 3895 24448 3959 24452
rect 3975 24508 4039 24512
rect 3975 24452 3979 24508
rect 3979 24452 4035 24508
rect 4035 24452 4039 24508
rect 3975 24448 4039 24452
rect 4055 24508 4119 24512
rect 4055 24452 4059 24508
rect 4059 24452 4115 24508
rect 4115 24452 4119 24508
rect 4055 24448 4119 24452
rect 9542 24508 9606 24512
rect 9542 24452 9546 24508
rect 9546 24452 9602 24508
rect 9602 24452 9606 24508
rect 9542 24448 9606 24452
rect 9622 24508 9686 24512
rect 9622 24452 9626 24508
rect 9626 24452 9682 24508
rect 9682 24452 9686 24508
rect 9622 24448 9686 24452
rect 9702 24508 9766 24512
rect 9702 24452 9706 24508
rect 9706 24452 9762 24508
rect 9762 24452 9766 24508
rect 9702 24448 9766 24452
rect 9782 24508 9846 24512
rect 9782 24452 9786 24508
rect 9786 24452 9842 24508
rect 9842 24452 9846 24508
rect 9782 24448 9846 24452
rect 15269 24508 15333 24512
rect 15269 24452 15273 24508
rect 15273 24452 15329 24508
rect 15329 24452 15333 24508
rect 15269 24448 15333 24452
rect 15349 24508 15413 24512
rect 15349 24452 15353 24508
rect 15353 24452 15409 24508
rect 15409 24452 15413 24508
rect 15349 24448 15413 24452
rect 15429 24508 15493 24512
rect 15429 24452 15433 24508
rect 15433 24452 15489 24508
rect 15489 24452 15493 24508
rect 15429 24448 15493 24452
rect 15509 24508 15573 24512
rect 15509 24452 15513 24508
rect 15513 24452 15569 24508
rect 15569 24452 15573 24508
rect 15509 24448 15573 24452
rect 20996 24508 21060 24512
rect 20996 24452 21000 24508
rect 21000 24452 21056 24508
rect 21056 24452 21060 24508
rect 20996 24448 21060 24452
rect 21076 24508 21140 24512
rect 21076 24452 21080 24508
rect 21080 24452 21136 24508
rect 21136 24452 21140 24508
rect 21076 24448 21140 24452
rect 21156 24508 21220 24512
rect 21156 24452 21160 24508
rect 21160 24452 21216 24508
rect 21216 24452 21220 24508
rect 21156 24448 21220 24452
rect 21236 24508 21300 24512
rect 21236 24452 21240 24508
rect 21240 24452 21296 24508
rect 21296 24452 21300 24508
rect 21236 24448 21300 24452
rect 4475 23964 4539 23968
rect 4475 23908 4479 23964
rect 4479 23908 4535 23964
rect 4535 23908 4539 23964
rect 4475 23904 4539 23908
rect 4555 23964 4619 23968
rect 4555 23908 4559 23964
rect 4559 23908 4615 23964
rect 4615 23908 4619 23964
rect 4555 23904 4619 23908
rect 4635 23964 4699 23968
rect 4635 23908 4639 23964
rect 4639 23908 4695 23964
rect 4695 23908 4699 23964
rect 4635 23904 4699 23908
rect 4715 23964 4779 23968
rect 4715 23908 4719 23964
rect 4719 23908 4775 23964
rect 4775 23908 4779 23964
rect 4715 23904 4779 23908
rect 10202 23964 10266 23968
rect 10202 23908 10206 23964
rect 10206 23908 10262 23964
rect 10262 23908 10266 23964
rect 10202 23904 10266 23908
rect 10282 23964 10346 23968
rect 10282 23908 10286 23964
rect 10286 23908 10342 23964
rect 10342 23908 10346 23964
rect 10282 23904 10346 23908
rect 10362 23964 10426 23968
rect 10362 23908 10366 23964
rect 10366 23908 10422 23964
rect 10422 23908 10426 23964
rect 10362 23904 10426 23908
rect 10442 23964 10506 23968
rect 10442 23908 10446 23964
rect 10446 23908 10502 23964
rect 10502 23908 10506 23964
rect 10442 23904 10506 23908
rect 15929 23964 15993 23968
rect 15929 23908 15933 23964
rect 15933 23908 15989 23964
rect 15989 23908 15993 23964
rect 15929 23904 15993 23908
rect 16009 23964 16073 23968
rect 16009 23908 16013 23964
rect 16013 23908 16069 23964
rect 16069 23908 16073 23964
rect 16009 23904 16073 23908
rect 16089 23964 16153 23968
rect 16089 23908 16093 23964
rect 16093 23908 16149 23964
rect 16149 23908 16153 23964
rect 16089 23904 16153 23908
rect 16169 23964 16233 23968
rect 16169 23908 16173 23964
rect 16173 23908 16229 23964
rect 16229 23908 16233 23964
rect 16169 23904 16233 23908
rect 21656 23964 21720 23968
rect 21656 23908 21660 23964
rect 21660 23908 21716 23964
rect 21716 23908 21720 23964
rect 21656 23904 21720 23908
rect 21736 23964 21800 23968
rect 21736 23908 21740 23964
rect 21740 23908 21796 23964
rect 21796 23908 21800 23964
rect 21736 23904 21800 23908
rect 21816 23964 21880 23968
rect 21816 23908 21820 23964
rect 21820 23908 21876 23964
rect 21876 23908 21880 23964
rect 21816 23904 21880 23908
rect 21896 23964 21960 23968
rect 21896 23908 21900 23964
rect 21900 23908 21956 23964
rect 21956 23908 21960 23964
rect 21896 23904 21960 23908
rect 3815 23420 3879 23424
rect 3815 23364 3819 23420
rect 3819 23364 3875 23420
rect 3875 23364 3879 23420
rect 3815 23360 3879 23364
rect 3895 23420 3959 23424
rect 3895 23364 3899 23420
rect 3899 23364 3955 23420
rect 3955 23364 3959 23420
rect 3895 23360 3959 23364
rect 3975 23420 4039 23424
rect 3975 23364 3979 23420
rect 3979 23364 4035 23420
rect 4035 23364 4039 23420
rect 3975 23360 4039 23364
rect 4055 23420 4119 23424
rect 4055 23364 4059 23420
rect 4059 23364 4115 23420
rect 4115 23364 4119 23420
rect 4055 23360 4119 23364
rect 9542 23420 9606 23424
rect 9542 23364 9546 23420
rect 9546 23364 9602 23420
rect 9602 23364 9606 23420
rect 9542 23360 9606 23364
rect 9622 23420 9686 23424
rect 9622 23364 9626 23420
rect 9626 23364 9682 23420
rect 9682 23364 9686 23420
rect 9622 23360 9686 23364
rect 9702 23420 9766 23424
rect 9702 23364 9706 23420
rect 9706 23364 9762 23420
rect 9762 23364 9766 23420
rect 9702 23360 9766 23364
rect 9782 23420 9846 23424
rect 9782 23364 9786 23420
rect 9786 23364 9842 23420
rect 9842 23364 9846 23420
rect 9782 23360 9846 23364
rect 15269 23420 15333 23424
rect 15269 23364 15273 23420
rect 15273 23364 15329 23420
rect 15329 23364 15333 23420
rect 15269 23360 15333 23364
rect 15349 23420 15413 23424
rect 15349 23364 15353 23420
rect 15353 23364 15409 23420
rect 15409 23364 15413 23420
rect 15349 23360 15413 23364
rect 15429 23420 15493 23424
rect 15429 23364 15433 23420
rect 15433 23364 15489 23420
rect 15489 23364 15493 23420
rect 15429 23360 15493 23364
rect 15509 23420 15573 23424
rect 15509 23364 15513 23420
rect 15513 23364 15569 23420
rect 15569 23364 15573 23420
rect 15509 23360 15573 23364
rect 20996 23420 21060 23424
rect 20996 23364 21000 23420
rect 21000 23364 21056 23420
rect 21056 23364 21060 23420
rect 20996 23360 21060 23364
rect 21076 23420 21140 23424
rect 21076 23364 21080 23420
rect 21080 23364 21136 23420
rect 21136 23364 21140 23420
rect 21076 23360 21140 23364
rect 21156 23420 21220 23424
rect 21156 23364 21160 23420
rect 21160 23364 21216 23420
rect 21216 23364 21220 23420
rect 21156 23360 21220 23364
rect 21236 23420 21300 23424
rect 21236 23364 21240 23420
rect 21240 23364 21296 23420
rect 21296 23364 21300 23420
rect 21236 23360 21300 23364
rect 4475 22876 4539 22880
rect 4475 22820 4479 22876
rect 4479 22820 4535 22876
rect 4535 22820 4539 22876
rect 4475 22816 4539 22820
rect 4555 22876 4619 22880
rect 4555 22820 4559 22876
rect 4559 22820 4615 22876
rect 4615 22820 4619 22876
rect 4555 22816 4619 22820
rect 4635 22876 4699 22880
rect 4635 22820 4639 22876
rect 4639 22820 4695 22876
rect 4695 22820 4699 22876
rect 4635 22816 4699 22820
rect 4715 22876 4779 22880
rect 4715 22820 4719 22876
rect 4719 22820 4775 22876
rect 4775 22820 4779 22876
rect 4715 22816 4779 22820
rect 10202 22876 10266 22880
rect 10202 22820 10206 22876
rect 10206 22820 10262 22876
rect 10262 22820 10266 22876
rect 10202 22816 10266 22820
rect 10282 22876 10346 22880
rect 10282 22820 10286 22876
rect 10286 22820 10342 22876
rect 10342 22820 10346 22876
rect 10282 22816 10346 22820
rect 10362 22876 10426 22880
rect 10362 22820 10366 22876
rect 10366 22820 10422 22876
rect 10422 22820 10426 22876
rect 10362 22816 10426 22820
rect 10442 22876 10506 22880
rect 10442 22820 10446 22876
rect 10446 22820 10502 22876
rect 10502 22820 10506 22876
rect 10442 22816 10506 22820
rect 15929 22876 15993 22880
rect 15929 22820 15933 22876
rect 15933 22820 15989 22876
rect 15989 22820 15993 22876
rect 15929 22816 15993 22820
rect 16009 22876 16073 22880
rect 16009 22820 16013 22876
rect 16013 22820 16069 22876
rect 16069 22820 16073 22876
rect 16009 22816 16073 22820
rect 16089 22876 16153 22880
rect 16089 22820 16093 22876
rect 16093 22820 16149 22876
rect 16149 22820 16153 22876
rect 16089 22816 16153 22820
rect 16169 22876 16233 22880
rect 16169 22820 16173 22876
rect 16173 22820 16229 22876
rect 16229 22820 16233 22876
rect 16169 22816 16233 22820
rect 21656 22876 21720 22880
rect 21656 22820 21660 22876
rect 21660 22820 21716 22876
rect 21716 22820 21720 22876
rect 21656 22816 21720 22820
rect 21736 22876 21800 22880
rect 21736 22820 21740 22876
rect 21740 22820 21796 22876
rect 21796 22820 21800 22876
rect 21736 22816 21800 22820
rect 21816 22876 21880 22880
rect 21816 22820 21820 22876
rect 21820 22820 21876 22876
rect 21876 22820 21880 22876
rect 21816 22816 21880 22820
rect 21896 22876 21960 22880
rect 21896 22820 21900 22876
rect 21900 22820 21956 22876
rect 21956 22820 21960 22876
rect 21896 22816 21960 22820
rect 3815 22332 3879 22336
rect 3815 22276 3819 22332
rect 3819 22276 3875 22332
rect 3875 22276 3879 22332
rect 3815 22272 3879 22276
rect 3895 22332 3959 22336
rect 3895 22276 3899 22332
rect 3899 22276 3955 22332
rect 3955 22276 3959 22332
rect 3895 22272 3959 22276
rect 3975 22332 4039 22336
rect 3975 22276 3979 22332
rect 3979 22276 4035 22332
rect 4035 22276 4039 22332
rect 3975 22272 4039 22276
rect 4055 22332 4119 22336
rect 4055 22276 4059 22332
rect 4059 22276 4115 22332
rect 4115 22276 4119 22332
rect 4055 22272 4119 22276
rect 9542 22332 9606 22336
rect 9542 22276 9546 22332
rect 9546 22276 9602 22332
rect 9602 22276 9606 22332
rect 9542 22272 9606 22276
rect 9622 22332 9686 22336
rect 9622 22276 9626 22332
rect 9626 22276 9682 22332
rect 9682 22276 9686 22332
rect 9622 22272 9686 22276
rect 9702 22332 9766 22336
rect 9702 22276 9706 22332
rect 9706 22276 9762 22332
rect 9762 22276 9766 22332
rect 9702 22272 9766 22276
rect 9782 22332 9846 22336
rect 9782 22276 9786 22332
rect 9786 22276 9842 22332
rect 9842 22276 9846 22332
rect 9782 22272 9846 22276
rect 15269 22332 15333 22336
rect 15269 22276 15273 22332
rect 15273 22276 15329 22332
rect 15329 22276 15333 22332
rect 15269 22272 15333 22276
rect 15349 22332 15413 22336
rect 15349 22276 15353 22332
rect 15353 22276 15409 22332
rect 15409 22276 15413 22332
rect 15349 22272 15413 22276
rect 15429 22332 15493 22336
rect 15429 22276 15433 22332
rect 15433 22276 15489 22332
rect 15489 22276 15493 22332
rect 15429 22272 15493 22276
rect 15509 22332 15573 22336
rect 15509 22276 15513 22332
rect 15513 22276 15569 22332
rect 15569 22276 15573 22332
rect 15509 22272 15573 22276
rect 20996 22332 21060 22336
rect 20996 22276 21000 22332
rect 21000 22276 21056 22332
rect 21056 22276 21060 22332
rect 20996 22272 21060 22276
rect 21076 22332 21140 22336
rect 21076 22276 21080 22332
rect 21080 22276 21136 22332
rect 21136 22276 21140 22332
rect 21076 22272 21140 22276
rect 21156 22332 21220 22336
rect 21156 22276 21160 22332
rect 21160 22276 21216 22332
rect 21216 22276 21220 22332
rect 21156 22272 21220 22276
rect 21236 22332 21300 22336
rect 21236 22276 21240 22332
rect 21240 22276 21296 22332
rect 21296 22276 21300 22332
rect 21236 22272 21300 22276
rect 4475 21788 4539 21792
rect 4475 21732 4479 21788
rect 4479 21732 4535 21788
rect 4535 21732 4539 21788
rect 4475 21728 4539 21732
rect 4555 21788 4619 21792
rect 4555 21732 4559 21788
rect 4559 21732 4615 21788
rect 4615 21732 4619 21788
rect 4555 21728 4619 21732
rect 4635 21788 4699 21792
rect 4635 21732 4639 21788
rect 4639 21732 4695 21788
rect 4695 21732 4699 21788
rect 4635 21728 4699 21732
rect 4715 21788 4779 21792
rect 4715 21732 4719 21788
rect 4719 21732 4775 21788
rect 4775 21732 4779 21788
rect 4715 21728 4779 21732
rect 10202 21788 10266 21792
rect 10202 21732 10206 21788
rect 10206 21732 10262 21788
rect 10262 21732 10266 21788
rect 10202 21728 10266 21732
rect 10282 21788 10346 21792
rect 10282 21732 10286 21788
rect 10286 21732 10342 21788
rect 10342 21732 10346 21788
rect 10282 21728 10346 21732
rect 10362 21788 10426 21792
rect 10362 21732 10366 21788
rect 10366 21732 10422 21788
rect 10422 21732 10426 21788
rect 10362 21728 10426 21732
rect 10442 21788 10506 21792
rect 10442 21732 10446 21788
rect 10446 21732 10502 21788
rect 10502 21732 10506 21788
rect 10442 21728 10506 21732
rect 15929 21788 15993 21792
rect 15929 21732 15933 21788
rect 15933 21732 15989 21788
rect 15989 21732 15993 21788
rect 15929 21728 15993 21732
rect 16009 21788 16073 21792
rect 16009 21732 16013 21788
rect 16013 21732 16069 21788
rect 16069 21732 16073 21788
rect 16009 21728 16073 21732
rect 16089 21788 16153 21792
rect 16089 21732 16093 21788
rect 16093 21732 16149 21788
rect 16149 21732 16153 21788
rect 16089 21728 16153 21732
rect 16169 21788 16233 21792
rect 16169 21732 16173 21788
rect 16173 21732 16229 21788
rect 16229 21732 16233 21788
rect 16169 21728 16233 21732
rect 21656 21788 21720 21792
rect 21656 21732 21660 21788
rect 21660 21732 21716 21788
rect 21716 21732 21720 21788
rect 21656 21728 21720 21732
rect 21736 21788 21800 21792
rect 21736 21732 21740 21788
rect 21740 21732 21796 21788
rect 21796 21732 21800 21788
rect 21736 21728 21800 21732
rect 21816 21788 21880 21792
rect 21816 21732 21820 21788
rect 21820 21732 21876 21788
rect 21876 21732 21880 21788
rect 21816 21728 21880 21732
rect 21896 21788 21960 21792
rect 21896 21732 21900 21788
rect 21900 21732 21956 21788
rect 21956 21732 21960 21788
rect 21896 21728 21960 21732
rect 3815 21244 3879 21248
rect 3815 21188 3819 21244
rect 3819 21188 3875 21244
rect 3875 21188 3879 21244
rect 3815 21184 3879 21188
rect 3895 21244 3959 21248
rect 3895 21188 3899 21244
rect 3899 21188 3955 21244
rect 3955 21188 3959 21244
rect 3895 21184 3959 21188
rect 3975 21244 4039 21248
rect 3975 21188 3979 21244
rect 3979 21188 4035 21244
rect 4035 21188 4039 21244
rect 3975 21184 4039 21188
rect 4055 21244 4119 21248
rect 4055 21188 4059 21244
rect 4059 21188 4115 21244
rect 4115 21188 4119 21244
rect 4055 21184 4119 21188
rect 9542 21244 9606 21248
rect 9542 21188 9546 21244
rect 9546 21188 9602 21244
rect 9602 21188 9606 21244
rect 9542 21184 9606 21188
rect 9622 21244 9686 21248
rect 9622 21188 9626 21244
rect 9626 21188 9682 21244
rect 9682 21188 9686 21244
rect 9622 21184 9686 21188
rect 9702 21244 9766 21248
rect 9702 21188 9706 21244
rect 9706 21188 9762 21244
rect 9762 21188 9766 21244
rect 9702 21184 9766 21188
rect 9782 21244 9846 21248
rect 9782 21188 9786 21244
rect 9786 21188 9842 21244
rect 9842 21188 9846 21244
rect 9782 21184 9846 21188
rect 15269 21244 15333 21248
rect 15269 21188 15273 21244
rect 15273 21188 15329 21244
rect 15329 21188 15333 21244
rect 15269 21184 15333 21188
rect 15349 21244 15413 21248
rect 15349 21188 15353 21244
rect 15353 21188 15409 21244
rect 15409 21188 15413 21244
rect 15349 21184 15413 21188
rect 15429 21244 15493 21248
rect 15429 21188 15433 21244
rect 15433 21188 15489 21244
rect 15489 21188 15493 21244
rect 15429 21184 15493 21188
rect 15509 21244 15573 21248
rect 15509 21188 15513 21244
rect 15513 21188 15569 21244
rect 15569 21188 15573 21244
rect 15509 21184 15573 21188
rect 20996 21244 21060 21248
rect 20996 21188 21000 21244
rect 21000 21188 21056 21244
rect 21056 21188 21060 21244
rect 20996 21184 21060 21188
rect 21076 21244 21140 21248
rect 21076 21188 21080 21244
rect 21080 21188 21136 21244
rect 21136 21188 21140 21244
rect 21076 21184 21140 21188
rect 21156 21244 21220 21248
rect 21156 21188 21160 21244
rect 21160 21188 21216 21244
rect 21216 21188 21220 21244
rect 21156 21184 21220 21188
rect 21236 21244 21300 21248
rect 21236 21188 21240 21244
rect 21240 21188 21296 21244
rect 21296 21188 21300 21244
rect 21236 21184 21300 21188
rect 4475 20700 4539 20704
rect 4475 20644 4479 20700
rect 4479 20644 4535 20700
rect 4535 20644 4539 20700
rect 4475 20640 4539 20644
rect 4555 20700 4619 20704
rect 4555 20644 4559 20700
rect 4559 20644 4615 20700
rect 4615 20644 4619 20700
rect 4555 20640 4619 20644
rect 4635 20700 4699 20704
rect 4635 20644 4639 20700
rect 4639 20644 4695 20700
rect 4695 20644 4699 20700
rect 4635 20640 4699 20644
rect 4715 20700 4779 20704
rect 4715 20644 4719 20700
rect 4719 20644 4775 20700
rect 4775 20644 4779 20700
rect 4715 20640 4779 20644
rect 10202 20700 10266 20704
rect 10202 20644 10206 20700
rect 10206 20644 10262 20700
rect 10262 20644 10266 20700
rect 10202 20640 10266 20644
rect 10282 20700 10346 20704
rect 10282 20644 10286 20700
rect 10286 20644 10342 20700
rect 10342 20644 10346 20700
rect 10282 20640 10346 20644
rect 10362 20700 10426 20704
rect 10362 20644 10366 20700
rect 10366 20644 10422 20700
rect 10422 20644 10426 20700
rect 10362 20640 10426 20644
rect 10442 20700 10506 20704
rect 10442 20644 10446 20700
rect 10446 20644 10502 20700
rect 10502 20644 10506 20700
rect 10442 20640 10506 20644
rect 15929 20700 15993 20704
rect 15929 20644 15933 20700
rect 15933 20644 15989 20700
rect 15989 20644 15993 20700
rect 15929 20640 15993 20644
rect 16009 20700 16073 20704
rect 16009 20644 16013 20700
rect 16013 20644 16069 20700
rect 16069 20644 16073 20700
rect 16009 20640 16073 20644
rect 16089 20700 16153 20704
rect 16089 20644 16093 20700
rect 16093 20644 16149 20700
rect 16149 20644 16153 20700
rect 16089 20640 16153 20644
rect 16169 20700 16233 20704
rect 16169 20644 16173 20700
rect 16173 20644 16229 20700
rect 16229 20644 16233 20700
rect 16169 20640 16233 20644
rect 21656 20700 21720 20704
rect 21656 20644 21660 20700
rect 21660 20644 21716 20700
rect 21716 20644 21720 20700
rect 21656 20640 21720 20644
rect 21736 20700 21800 20704
rect 21736 20644 21740 20700
rect 21740 20644 21796 20700
rect 21796 20644 21800 20700
rect 21736 20640 21800 20644
rect 21816 20700 21880 20704
rect 21816 20644 21820 20700
rect 21820 20644 21876 20700
rect 21876 20644 21880 20700
rect 21816 20640 21880 20644
rect 21896 20700 21960 20704
rect 21896 20644 21900 20700
rect 21900 20644 21956 20700
rect 21956 20644 21960 20700
rect 21896 20640 21960 20644
rect 3815 20156 3879 20160
rect 3815 20100 3819 20156
rect 3819 20100 3875 20156
rect 3875 20100 3879 20156
rect 3815 20096 3879 20100
rect 3895 20156 3959 20160
rect 3895 20100 3899 20156
rect 3899 20100 3955 20156
rect 3955 20100 3959 20156
rect 3895 20096 3959 20100
rect 3975 20156 4039 20160
rect 3975 20100 3979 20156
rect 3979 20100 4035 20156
rect 4035 20100 4039 20156
rect 3975 20096 4039 20100
rect 4055 20156 4119 20160
rect 4055 20100 4059 20156
rect 4059 20100 4115 20156
rect 4115 20100 4119 20156
rect 4055 20096 4119 20100
rect 9542 20156 9606 20160
rect 9542 20100 9546 20156
rect 9546 20100 9602 20156
rect 9602 20100 9606 20156
rect 9542 20096 9606 20100
rect 9622 20156 9686 20160
rect 9622 20100 9626 20156
rect 9626 20100 9682 20156
rect 9682 20100 9686 20156
rect 9622 20096 9686 20100
rect 9702 20156 9766 20160
rect 9702 20100 9706 20156
rect 9706 20100 9762 20156
rect 9762 20100 9766 20156
rect 9702 20096 9766 20100
rect 9782 20156 9846 20160
rect 9782 20100 9786 20156
rect 9786 20100 9842 20156
rect 9842 20100 9846 20156
rect 9782 20096 9846 20100
rect 15269 20156 15333 20160
rect 15269 20100 15273 20156
rect 15273 20100 15329 20156
rect 15329 20100 15333 20156
rect 15269 20096 15333 20100
rect 15349 20156 15413 20160
rect 15349 20100 15353 20156
rect 15353 20100 15409 20156
rect 15409 20100 15413 20156
rect 15349 20096 15413 20100
rect 15429 20156 15493 20160
rect 15429 20100 15433 20156
rect 15433 20100 15489 20156
rect 15489 20100 15493 20156
rect 15429 20096 15493 20100
rect 15509 20156 15573 20160
rect 15509 20100 15513 20156
rect 15513 20100 15569 20156
rect 15569 20100 15573 20156
rect 15509 20096 15573 20100
rect 20996 20156 21060 20160
rect 20996 20100 21000 20156
rect 21000 20100 21056 20156
rect 21056 20100 21060 20156
rect 20996 20096 21060 20100
rect 21076 20156 21140 20160
rect 21076 20100 21080 20156
rect 21080 20100 21136 20156
rect 21136 20100 21140 20156
rect 21076 20096 21140 20100
rect 21156 20156 21220 20160
rect 21156 20100 21160 20156
rect 21160 20100 21216 20156
rect 21216 20100 21220 20156
rect 21156 20096 21220 20100
rect 21236 20156 21300 20160
rect 21236 20100 21240 20156
rect 21240 20100 21296 20156
rect 21296 20100 21300 20156
rect 21236 20096 21300 20100
rect 4475 19612 4539 19616
rect 4475 19556 4479 19612
rect 4479 19556 4535 19612
rect 4535 19556 4539 19612
rect 4475 19552 4539 19556
rect 4555 19612 4619 19616
rect 4555 19556 4559 19612
rect 4559 19556 4615 19612
rect 4615 19556 4619 19612
rect 4555 19552 4619 19556
rect 4635 19612 4699 19616
rect 4635 19556 4639 19612
rect 4639 19556 4695 19612
rect 4695 19556 4699 19612
rect 4635 19552 4699 19556
rect 4715 19612 4779 19616
rect 4715 19556 4719 19612
rect 4719 19556 4775 19612
rect 4775 19556 4779 19612
rect 4715 19552 4779 19556
rect 10202 19612 10266 19616
rect 10202 19556 10206 19612
rect 10206 19556 10262 19612
rect 10262 19556 10266 19612
rect 10202 19552 10266 19556
rect 10282 19612 10346 19616
rect 10282 19556 10286 19612
rect 10286 19556 10342 19612
rect 10342 19556 10346 19612
rect 10282 19552 10346 19556
rect 10362 19612 10426 19616
rect 10362 19556 10366 19612
rect 10366 19556 10422 19612
rect 10422 19556 10426 19612
rect 10362 19552 10426 19556
rect 10442 19612 10506 19616
rect 10442 19556 10446 19612
rect 10446 19556 10502 19612
rect 10502 19556 10506 19612
rect 10442 19552 10506 19556
rect 15929 19612 15993 19616
rect 15929 19556 15933 19612
rect 15933 19556 15989 19612
rect 15989 19556 15993 19612
rect 15929 19552 15993 19556
rect 16009 19612 16073 19616
rect 16009 19556 16013 19612
rect 16013 19556 16069 19612
rect 16069 19556 16073 19612
rect 16009 19552 16073 19556
rect 16089 19612 16153 19616
rect 16089 19556 16093 19612
rect 16093 19556 16149 19612
rect 16149 19556 16153 19612
rect 16089 19552 16153 19556
rect 16169 19612 16233 19616
rect 16169 19556 16173 19612
rect 16173 19556 16229 19612
rect 16229 19556 16233 19612
rect 16169 19552 16233 19556
rect 21656 19612 21720 19616
rect 21656 19556 21660 19612
rect 21660 19556 21716 19612
rect 21716 19556 21720 19612
rect 21656 19552 21720 19556
rect 21736 19612 21800 19616
rect 21736 19556 21740 19612
rect 21740 19556 21796 19612
rect 21796 19556 21800 19612
rect 21736 19552 21800 19556
rect 21816 19612 21880 19616
rect 21816 19556 21820 19612
rect 21820 19556 21876 19612
rect 21876 19556 21880 19612
rect 21816 19552 21880 19556
rect 21896 19612 21960 19616
rect 21896 19556 21900 19612
rect 21900 19556 21956 19612
rect 21956 19556 21960 19612
rect 21896 19552 21960 19556
rect 3815 19068 3879 19072
rect 3815 19012 3819 19068
rect 3819 19012 3875 19068
rect 3875 19012 3879 19068
rect 3815 19008 3879 19012
rect 3895 19068 3959 19072
rect 3895 19012 3899 19068
rect 3899 19012 3955 19068
rect 3955 19012 3959 19068
rect 3895 19008 3959 19012
rect 3975 19068 4039 19072
rect 3975 19012 3979 19068
rect 3979 19012 4035 19068
rect 4035 19012 4039 19068
rect 3975 19008 4039 19012
rect 4055 19068 4119 19072
rect 4055 19012 4059 19068
rect 4059 19012 4115 19068
rect 4115 19012 4119 19068
rect 4055 19008 4119 19012
rect 9542 19068 9606 19072
rect 9542 19012 9546 19068
rect 9546 19012 9602 19068
rect 9602 19012 9606 19068
rect 9542 19008 9606 19012
rect 9622 19068 9686 19072
rect 9622 19012 9626 19068
rect 9626 19012 9682 19068
rect 9682 19012 9686 19068
rect 9622 19008 9686 19012
rect 9702 19068 9766 19072
rect 9702 19012 9706 19068
rect 9706 19012 9762 19068
rect 9762 19012 9766 19068
rect 9702 19008 9766 19012
rect 9782 19068 9846 19072
rect 9782 19012 9786 19068
rect 9786 19012 9842 19068
rect 9842 19012 9846 19068
rect 9782 19008 9846 19012
rect 15269 19068 15333 19072
rect 15269 19012 15273 19068
rect 15273 19012 15329 19068
rect 15329 19012 15333 19068
rect 15269 19008 15333 19012
rect 15349 19068 15413 19072
rect 15349 19012 15353 19068
rect 15353 19012 15409 19068
rect 15409 19012 15413 19068
rect 15349 19008 15413 19012
rect 15429 19068 15493 19072
rect 15429 19012 15433 19068
rect 15433 19012 15489 19068
rect 15489 19012 15493 19068
rect 15429 19008 15493 19012
rect 15509 19068 15573 19072
rect 15509 19012 15513 19068
rect 15513 19012 15569 19068
rect 15569 19012 15573 19068
rect 15509 19008 15573 19012
rect 20996 19068 21060 19072
rect 20996 19012 21000 19068
rect 21000 19012 21056 19068
rect 21056 19012 21060 19068
rect 20996 19008 21060 19012
rect 21076 19068 21140 19072
rect 21076 19012 21080 19068
rect 21080 19012 21136 19068
rect 21136 19012 21140 19068
rect 21076 19008 21140 19012
rect 21156 19068 21220 19072
rect 21156 19012 21160 19068
rect 21160 19012 21216 19068
rect 21216 19012 21220 19068
rect 21156 19008 21220 19012
rect 21236 19068 21300 19072
rect 21236 19012 21240 19068
rect 21240 19012 21296 19068
rect 21296 19012 21300 19068
rect 21236 19008 21300 19012
rect 4475 18524 4539 18528
rect 4475 18468 4479 18524
rect 4479 18468 4535 18524
rect 4535 18468 4539 18524
rect 4475 18464 4539 18468
rect 4555 18524 4619 18528
rect 4555 18468 4559 18524
rect 4559 18468 4615 18524
rect 4615 18468 4619 18524
rect 4555 18464 4619 18468
rect 4635 18524 4699 18528
rect 4635 18468 4639 18524
rect 4639 18468 4695 18524
rect 4695 18468 4699 18524
rect 4635 18464 4699 18468
rect 4715 18524 4779 18528
rect 4715 18468 4719 18524
rect 4719 18468 4775 18524
rect 4775 18468 4779 18524
rect 4715 18464 4779 18468
rect 10202 18524 10266 18528
rect 10202 18468 10206 18524
rect 10206 18468 10262 18524
rect 10262 18468 10266 18524
rect 10202 18464 10266 18468
rect 10282 18524 10346 18528
rect 10282 18468 10286 18524
rect 10286 18468 10342 18524
rect 10342 18468 10346 18524
rect 10282 18464 10346 18468
rect 10362 18524 10426 18528
rect 10362 18468 10366 18524
rect 10366 18468 10422 18524
rect 10422 18468 10426 18524
rect 10362 18464 10426 18468
rect 10442 18524 10506 18528
rect 10442 18468 10446 18524
rect 10446 18468 10502 18524
rect 10502 18468 10506 18524
rect 10442 18464 10506 18468
rect 15929 18524 15993 18528
rect 15929 18468 15933 18524
rect 15933 18468 15989 18524
rect 15989 18468 15993 18524
rect 15929 18464 15993 18468
rect 16009 18524 16073 18528
rect 16009 18468 16013 18524
rect 16013 18468 16069 18524
rect 16069 18468 16073 18524
rect 16009 18464 16073 18468
rect 16089 18524 16153 18528
rect 16089 18468 16093 18524
rect 16093 18468 16149 18524
rect 16149 18468 16153 18524
rect 16089 18464 16153 18468
rect 16169 18524 16233 18528
rect 16169 18468 16173 18524
rect 16173 18468 16229 18524
rect 16229 18468 16233 18524
rect 16169 18464 16233 18468
rect 21656 18524 21720 18528
rect 21656 18468 21660 18524
rect 21660 18468 21716 18524
rect 21716 18468 21720 18524
rect 21656 18464 21720 18468
rect 21736 18524 21800 18528
rect 21736 18468 21740 18524
rect 21740 18468 21796 18524
rect 21796 18468 21800 18524
rect 21736 18464 21800 18468
rect 21816 18524 21880 18528
rect 21816 18468 21820 18524
rect 21820 18468 21876 18524
rect 21876 18468 21880 18524
rect 21816 18464 21880 18468
rect 21896 18524 21960 18528
rect 21896 18468 21900 18524
rect 21900 18468 21956 18524
rect 21956 18468 21960 18524
rect 21896 18464 21960 18468
rect 3815 17980 3879 17984
rect 3815 17924 3819 17980
rect 3819 17924 3875 17980
rect 3875 17924 3879 17980
rect 3815 17920 3879 17924
rect 3895 17980 3959 17984
rect 3895 17924 3899 17980
rect 3899 17924 3955 17980
rect 3955 17924 3959 17980
rect 3895 17920 3959 17924
rect 3975 17980 4039 17984
rect 3975 17924 3979 17980
rect 3979 17924 4035 17980
rect 4035 17924 4039 17980
rect 3975 17920 4039 17924
rect 4055 17980 4119 17984
rect 4055 17924 4059 17980
rect 4059 17924 4115 17980
rect 4115 17924 4119 17980
rect 4055 17920 4119 17924
rect 9542 17980 9606 17984
rect 9542 17924 9546 17980
rect 9546 17924 9602 17980
rect 9602 17924 9606 17980
rect 9542 17920 9606 17924
rect 9622 17980 9686 17984
rect 9622 17924 9626 17980
rect 9626 17924 9682 17980
rect 9682 17924 9686 17980
rect 9622 17920 9686 17924
rect 9702 17980 9766 17984
rect 9702 17924 9706 17980
rect 9706 17924 9762 17980
rect 9762 17924 9766 17980
rect 9702 17920 9766 17924
rect 9782 17980 9846 17984
rect 9782 17924 9786 17980
rect 9786 17924 9842 17980
rect 9842 17924 9846 17980
rect 9782 17920 9846 17924
rect 15269 17980 15333 17984
rect 15269 17924 15273 17980
rect 15273 17924 15329 17980
rect 15329 17924 15333 17980
rect 15269 17920 15333 17924
rect 15349 17980 15413 17984
rect 15349 17924 15353 17980
rect 15353 17924 15409 17980
rect 15409 17924 15413 17980
rect 15349 17920 15413 17924
rect 15429 17980 15493 17984
rect 15429 17924 15433 17980
rect 15433 17924 15489 17980
rect 15489 17924 15493 17980
rect 15429 17920 15493 17924
rect 15509 17980 15573 17984
rect 15509 17924 15513 17980
rect 15513 17924 15569 17980
rect 15569 17924 15573 17980
rect 15509 17920 15573 17924
rect 20996 17980 21060 17984
rect 20996 17924 21000 17980
rect 21000 17924 21056 17980
rect 21056 17924 21060 17980
rect 20996 17920 21060 17924
rect 21076 17980 21140 17984
rect 21076 17924 21080 17980
rect 21080 17924 21136 17980
rect 21136 17924 21140 17980
rect 21076 17920 21140 17924
rect 21156 17980 21220 17984
rect 21156 17924 21160 17980
rect 21160 17924 21216 17980
rect 21216 17924 21220 17980
rect 21156 17920 21220 17924
rect 21236 17980 21300 17984
rect 21236 17924 21240 17980
rect 21240 17924 21296 17980
rect 21296 17924 21300 17980
rect 21236 17920 21300 17924
rect 4475 17436 4539 17440
rect 4475 17380 4479 17436
rect 4479 17380 4535 17436
rect 4535 17380 4539 17436
rect 4475 17376 4539 17380
rect 4555 17436 4619 17440
rect 4555 17380 4559 17436
rect 4559 17380 4615 17436
rect 4615 17380 4619 17436
rect 4555 17376 4619 17380
rect 4635 17436 4699 17440
rect 4635 17380 4639 17436
rect 4639 17380 4695 17436
rect 4695 17380 4699 17436
rect 4635 17376 4699 17380
rect 4715 17436 4779 17440
rect 4715 17380 4719 17436
rect 4719 17380 4775 17436
rect 4775 17380 4779 17436
rect 4715 17376 4779 17380
rect 10202 17436 10266 17440
rect 10202 17380 10206 17436
rect 10206 17380 10262 17436
rect 10262 17380 10266 17436
rect 10202 17376 10266 17380
rect 10282 17436 10346 17440
rect 10282 17380 10286 17436
rect 10286 17380 10342 17436
rect 10342 17380 10346 17436
rect 10282 17376 10346 17380
rect 10362 17436 10426 17440
rect 10362 17380 10366 17436
rect 10366 17380 10422 17436
rect 10422 17380 10426 17436
rect 10362 17376 10426 17380
rect 10442 17436 10506 17440
rect 10442 17380 10446 17436
rect 10446 17380 10502 17436
rect 10502 17380 10506 17436
rect 10442 17376 10506 17380
rect 15929 17436 15993 17440
rect 15929 17380 15933 17436
rect 15933 17380 15989 17436
rect 15989 17380 15993 17436
rect 15929 17376 15993 17380
rect 16009 17436 16073 17440
rect 16009 17380 16013 17436
rect 16013 17380 16069 17436
rect 16069 17380 16073 17436
rect 16009 17376 16073 17380
rect 16089 17436 16153 17440
rect 16089 17380 16093 17436
rect 16093 17380 16149 17436
rect 16149 17380 16153 17436
rect 16089 17376 16153 17380
rect 16169 17436 16233 17440
rect 16169 17380 16173 17436
rect 16173 17380 16229 17436
rect 16229 17380 16233 17436
rect 16169 17376 16233 17380
rect 21656 17436 21720 17440
rect 21656 17380 21660 17436
rect 21660 17380 21716 17436
rect 21716 17380 21720 17436
rect 21656 17376 21720 17380
rect 21736 17436 21800 17440
rect 21736 17380 21740 17436
rect 21740 17380 21796 17436
rect 21796 17380 21800 17436
rect 21736 17376 21800 17380
rect 21816 17436 21880 17440
rect 21816 17380 21820 17436
rect 21820 17380 21876 17436
rect 21876 17380 21880 17436
rect 21816 17376 21880 17380
rect 21896 17436 21960 17440
rect 21896 17380 21900 17436
rect 21900 17380 21956 17436
rect 21956 17380 21960 17436
rect 21896 17376 21960 17380
rect 3815 16892 3879 16896
rect 3815 16836 3819 16892
rect 3819 16836 3875 16892
rect 3875 16836 3879 16892
rect 3815 16832 3879 16836
rect 3895 16892 3959 16896
rect 3895 16836 3899 16892
rect 3899 16836 3955 16892
rect 3955 16836 3959 16892
rect 3895 16832 3959 16836
rect 3975 16892 4039 16896
rect 3975 16836 3979 16892
rect 3979 16836 4035 16892
rect 4035 16836 4039 16892
rect 3975 16832 4039 16836
rect 4055 16892 4119 16896
rect 4055 16836 4059 16892
rect 4059 16836 4115 16892
rect 4115 16836 4119 16892
rect 4055 16832 4119 16836
rect 9542 16892 9606 16896
rect 9542 16836 9546 16892
rect 9546 16836 9602 16892
rect 9602 16836 9606 16892
rect 9542 16832 9606 16836
rect 9622 16892 9686 16896
rect 9622 16836 9626 16892
rect 9626 16836 9682 16892
rect 9682 16836 9686 16892
rect 9622 16832 9686 16836
rect 9702 16892 9766 16896
rect 9702 16836 9706 16892
rect 9706 16836 9762 16892
rect 9762 16836 9766 16892
rect 9702 16832 9766 16836
rect 9782 16892 9846 16896
rect 9782 16836 9786 16892
rect 9786 16836 9842 16892
rect 9842 16836 9846 16892
rect 9782 16832 9846 16836
rect 15269 16892 15333 16896
rect 15269 16836 15273 16892
rect 15273 16836 15329 16892
rect 15329 16836 15333 16892
rect 15269 16832 15333 16836
rect 15349 16892 15413 16896
rect 15349 16836 15353 16892
rect 15353 16836 15409 16892
rect 15409 16836 15413 16892
rect 15349 16832 15413 16836
rect 15429 16892 15493 16896
rect 15429 16836 15433 16892
rect 15433 16836 15489 16892
rect 15489 16836 15493 16892
rect 15429 16832 15493 16836
rect 15509 16892 15573 16896
rect 15509 16836 15513 16892
rect 15513 16836 15569 16892
rect 15569 16836 15573 16892
rect 15509 16832 15573 16836
rect 20996 16892 21060 16896
rect 20996 16836 21000 16892
rect 21000 16836 21056 16892
rect 21056 16836 21060 16892
rect 20996 16832 21060 16836
rect 21076 16892 21140 16896
rect 21076 16836 21080 16892
rect 21080 16836 21136 16892
rect 21136 16836 21140 16892
rect 21076 16832 21140 16836
rect 21156 16892 21220 16896
rect 21156 16836 21160 16892
rect 21160 16836 21216 16892
rect 21216 16836 21220 16892
rect 21156 16832 21220 16836
rect 21236 16892 21300 16896
rect 21236 16836 21240 16892
rect 21240 16836 21296 16892
rect 21296 16836 21300 16892
rect 21236 16832 21300 16836
rect 4475 16348 4539 16352
rect 4475 16292 4479 16348
rect 4479 16292 4535 16348
rect 4535 16292 4539 16348
rect 4475 16288 4539 16292
rect 4555 16348 4619 16352
rect 4555 16292 4559 16348
rect 4559 16292 4615 16348
rect 4615 16292 4619 16348
rect 4555 16288 4619 16292
rect 4635 16348 4699 16352
rect 4635 16292 4639 16348
rect 4639 16292 4695 16348
rect 4695 16292 4699 16348
rect 4635 16288 4699 16292
rect 4715 16348 4779 16352
rect 4715 16292 4719 16348
rect 4719 16292 4775 16348
rect 4775 16292 4779 16348
rect 4715 16288 4779 16292
rect 10202 16348 10266 16352
rect 10202 16292 10206 16348
rect 10206 16292 10262 16348
rect 10262 16292 10266 16348
rect 10202 16288 10266 16292
rect 10282 16348 10346 16352
rect 10282 16292 10286 16348
rect 10286 16292 10342 16348
rect 10342 16292 10346 16348
rect 10282 16288 10346 16292
rect 10362 16348 10426 16352
rect 10362 16292 10366 16348
rect 10366 16292 10422 16348
rect 10422 16292 10426 16348
rect 10362 16288 10426 16292
rect 10442 16348 10506 16352
rect 10442 16292 10446 16348
rect 10446 16292 10502 16348
rect 10502 16292 10506 16348
rect 10442 16288 10506 16292
rect 15929 16348 15993 16352
rect 15929 16292 15933 16348
rect 15933 16292 15989 16348
rect 15989 16292 15993 16348
rect 15929 16288 15993 16292
rect 16009 16348 16073 16352
rect 16009 16292 16013 16348
rect 16013 16292 16069 16348
rect 16069 16292 16073 16348
rect 16009 16288 16073 16292
rect 16089 16348 16153 16352
rect 16089 16292 16093 16348
rect 16093 16292 16149 16348
rect 16149 16292 16153 16348
rect 16089 16288 16153 16292
rect 16169 16348 16233 16352
rect 16169 16292 16173 16348
rect 16173 16292 16229 16348
rect 16229 16292 16233 16348
rect 16169 16288 16233 16292
rect 21656 16348 21720 16352
rect 21656 16292 21660 16348
rect 21660 16292 21716 16348
rect 21716 16292 21720 16348
rect 21656 16288 21720 16292
rect 21736 16348 21800 16352
rect 21736 16292 21740 16348
rect 21740 16292 21796 16348
rect 21796 16292 21800 16348
rect 21736 16288 21800 16292
rect 21816 16348 21880 16352
rect 21816 16292 21820 16348
rect 21820 16292 21876 16348
rect 21876 16292 21880 16348
rect 21816 16288 21880 16292
rect 21896 16348 21960 16352
rect 21896 16292 21900 16348
rect 21900 16292 21956 16348
rect 21956 16292 21960 16348
rect 21896 16288 21960 16292
rect 3815 15804 3879 15808
rect 3815 15748 3819 15804
rect 3819 15748 3875 15804
rect 3875 15748 3879 15804
rect 3815 15744 3879 15748
rect 3895 15804 3959 15808
rect 3895 15748 3899 15804
rect 3899 15748 3955 15804
rect 3955 15748 3959 15804
rect 3895 15744 3959 15748
rect 3975 15804 4039 15808
rect 3975 15748 3979 15804
rect 3979 15748 4035 15804
rect 4035 15748 4039 15804
rect 3975 15744 4039 15748
rect 4055 15804 4119 15808
rect 4055 15748 4059 15804
rect 4059 15748 4115 15804
rect 4115 15748 4119 15804
rect 4055 15744 4119 15748
rect 9542 15804 9606 15808
rect 9542 15748 9546 15804
rect 9546 15748 9602 15804
rect 9602 15748 9606 15804
rect 9542 15744 9606 15748
rect 9622 15804 9686 15808
rect 9622 15748 9626 15804
rect 9626 15748 9682 15804
rect 9682 15748 9686 15804
rect 9622 15744 9686 15748
rect 9702 15804 9766 15808
rect 9702 15748 9706 15804
rect 9706 15748 9762 15804
rect 9762 15748 9766 15804
rect 9702 15744 9766 15748
rect 9782 15804 9846 15808
rect 9782 15748 9786 15804
rect 9786 15748 9842 15804
rect 9842 15748 9846 15804
rect 9782 15744 9846 15748
rect 15269 15804 15333 15808
rect 15269 15748 15273 15804
rect 15273 15748 15329 15804
rect 15329 15748 15333 15804
rect 15269 15744 15333 15748
rect 15349 15804 15413 15808
rect 15349 15748 15353 15804
rect 15353 15748 15409 15804
rect 15409 15748 15413 15804
rect 15349 15744 15413 15748
rect 15429 15804 15493 15808
rect 15429 15748 15433 15804
rect 15433 15748 15489 15804
rect 15489 15748 15493 15804
rect 15429 15744 15493 15748
rect 15509 15804 15573 15808
rect 15509 15748 15513 15804
rect 15513 15748 15569 15804
rect 15569 15748 15573 15804
rect 15509 15744 15573 15748
rect 20996 15804 21060 15808
rect 20996 15748 21000 15804
rect 21000 15748 21056 15804
rect 21056 15748 21060 15804
rect 20996 15744 21060 15748
rect 21076 15804 21140 15808
rect 21076 15748 21080 15804
rect 21080 15748 21136 15804
rect 21136 15748 21140 15804
rect 21076 15744 21140 15748
rect 21156 15804 21220 15808
rect 21156 15748 21160 15804
rect 21160 15748 21216 15804
rect 21216 15748 21220 15804
rect 21156 15744 21220 15748
rect 21236 15804 21300 15808
rect 21236 15748 21240 15804
rect 21240 15748 21296 15804
rect 21296 15748 21300 15804
rect 21236 15744 21300 15748
rect 4475 15260 4539 15264
rect 4475 15204 4479 15260
rect 4479 15204 4535 15260
rect 4535 15204 4539 15260
rect 4475 15200 4539 15204
rect 4555 15260 4619 15264
rect 4555 15204 4559 15260
rect 4559 15204 4615 15260
rect 4615 15204 4619 15260
rect 4555 15200 4619 15204
rect 4635 15260 4699 15264
rect 4635 15204 4639 15260
rect 4639 15204 4695 15260
rect 4695 15204 4699 15260
rect 4635 15200 4699 15204
rect 4715 15260 4779 15264
rect 4715 15204 4719 15260
rect 4719 15204 4775 15260
rect 4775 15204 4779 15260
rect 4715 15200 4779 15204
rect 10202 15260 10266 15264
rect 10202 15204 10206 15260
rect 10206 15204 10262 15260
rect 10262 15204 10266 15260
rect 10202 15200 10266 15204
rect 10282 15260 10346 15264
rect 10282 15204 10286 15260
rect 10286 15204 10342 15260
rect 10342 15204 10346 15260
rect 10282 15200 10346 15204
rect 10362 15260 10426 15264
rect 10362 15204 10366 15260
rect 10366 15204 10422 15260
rect 10422 15204 10426 15260
rect 10362 15200 10426 15204
rect 10442 15260 10506 15264
rect 10442 15204 10446 15260
rect 10446 15204 10502 15260
rect 10502 15204 10506 15260
rect 10442 15200 10506 15204
rect 15929 15260 15993 15264
rect 15929 15204 15933 15260
rect 15933 15204 15989 15260
rect 15989 15204 15993 15260
rect 15929 15200 15993 15204
rect 16009 15260 16073 15264
rect 16009 15204 16013 15260
rect 16013 15204 16069 15260
rect 16069 15204 16073 15260
rect 16009 15200 16073 15204
rect 16089 15260 16153 15264
rect 16089 15204 16093 15260
rect 16093 15204 16149 15260
rect 16149 15204 16153 15260
rect 16089 15200 16153 15204
rect 16169 15260 16233 15264
rect 16169 15204 16173 15260
rect 16173 15204 16229 15260
rect 16229 15204 16233 15260
rect 16169 15200 16233 15204
rect 21656 15260 21720 15264
rect 21656 15204 21660 15260
rect 21660 15204 21716 15260
rect 21716 15204 21720 15260
rect 21656 15200 21720 15204
rect 21736 15260 21800 15264
rect 21736 15204 21740 15260
rect 21740 15204 21796 15260
rect 21796 15204 21800 15260
rect 21736 15200 21800 15204
rect 21816 15260 21880 15264
rect 21816 15204 21820 15260
rect 21820 15204 21876 15260
rect 21876 15204 21880 15260
rect 21816 15200 21880 15204
rect 21896 15260 21960 15264
rect 21896 15204 21900 15260
rect 21900 15204 21956 15260
rect 21956 15204 21960 15260
rect 21896 15200 21960 15204
rect 3815 14716 3879 14720
rect 3815 14660 3819 14716
rect 3819 14660 3875 14716
rect 3875 14660 3879 14716
rect 3815 14656 3879 14660
rect 3895 14716 3959 14720
rect 3895 14660 3899 14716
rect 3899 14660 3955 14716
rect 3955 14660 3959 14716
rect 3895 14656 3959 14660
rect 3975 14716 4039 14720
rect 3975 14660 3979 14716
rect 3979 14660 4035 14716
rect 4035 14660 4039 14716
rect 3975 14656 4039 14660
rect 4055 14716 4119 14720
rect 4055 14660 4059 14716
rect 4059 14660 4115 14716
rect 4115 14660 4119 14716
rect 4055 14656 4119 14660
rect 9542 14716 9606 14720
rect 9542 14660 9546 14716
rect 9546 14660 9602 14716
rect 9602 14660 9606 14716
rect 9542 14656 9606 14660
rect 9622 14716 9686 14720
rect 9622 14660 9626 14716
rect 9626 14660 9682 14716
rect 9682 14660 9686 14716
rect 9622 14656 9686 14660
rect 9702 14716 9766 14720
rect 9702 14660 9706 14716
rect 9706 14660 9762 14716
rect 9762 14660 9766 14716
rect 9702 14656 9766 14660
rect 9782 14716 9846 14720
rect 9782 14660 9786 14716
rect 9786 14660 9842 14716
rect 9842 14660 9846 14716
rect 9782 14656 9846 14660
rect 15269 14716 15333 14720
rect 15269 14660 15273 14716
rect 15273 14660 15329 14716
rect 15329 14660 15333 14716
rect 15269 14656 15333 14660
rect 15349 14716 15413 14720
rect 15349 14660 15353 14716
rect 15353 14660 15409 14716
rect 15409 14660 15413 14716
rect 15349 14656 15413 14660
rect 15429 14716 15493 14720
rect 15429 14660 15433 14716
rect 15433 14660 15489 14716
rect 15489 14660 15493 14716
rect 15429 14656 15493 14660
rect 15509 14716 15573 14720
rect 15509 14660 15513 14716
rect 15513 14660 15569 14716
rect 15569 14660 15573 14716
rect 15509 14656 15573 14660
rect 20996 14716 21060 14720
rect 20996 14660 21000 14716
rect 21000 14660 21056 14716
rect 21056 14660 21060 14716
rect 20996 14656 21060 14660
rect 21076 14716 21140 14720
rect 21076 14660 21080 14716
rect 21080 14660 21136 14716
rect 21136 14660 21140 14716
rect 21076 14656 21140 14660
rect 21156 14716 21220 14720
rect 21156 14660 21160 14716
rect 21160 14660 21216 14716
rect 21216 14660 21220 14716
rect 21156 14656 21220 14660
rect 21236 14716 21300 14720
rect 21236 14660 21240 14716
rect 21240 14660 21296 14716
rect 21296 14660 21300 14716
rect 21236 14656 21300 14660
rect 4475 14172 4539 14176
rect 4475 14116 4479 14172
rect 4479 14116 4535 14172
rect 4535 14116 4539 14172
rect 4475 14112 4539 14116
rect 4555 14172 4619 14176
rect 4555 14116 4559 14172
rect 4559 14116 4615 14172
rect 4615 14116 4619 14172
rect 4555 14112 4619 14116
rect 4635 14172 4699 14176
rect 4635 14116 4639 14172
rect 4639 14116 4695 14172
rect 4695 14116 4699 14172
rect 4635 14112 4699 14116
rect 4715 14172 4779 14176
rect 4715 14116 4719 14172
rect 4719 14116 4775 14172
rect 4775 14116 4779 14172
rect 4715 14112 4779 14116
rect 10202 14172 10266 14176
rect 10202 14116 10206 14172
rect 10206 14116 10262 14172
rect 10262 14116 10266 14172
rect 10202 14112 10266 14116
rect 10282 14172 10346 14176
rect 10282 14116 10286 14172
rect 10286 14116 10342 14172
rect 10342 14116 10346 14172
rect 10282 14112 10346 14116
rect 10362 14172 10426 14176
rect 10362 14116 10366 14172
rect 10366 14116 10422 14172
rect 10422 14116 10426 14172
rect 10362 14112 10426 14116
rect 10442 14172 10506 14176
rect 10442 14116 10446 14172
rect 10446 14116 10502 14172
rect 10502 14116 10506 14172
rect 10442 14112 10506 14116
rect 15929 14172 15993 14176
rect 15929 14116 15933 14172
rect 15933 14116 15989 14172
rect 15989 14116 15993 14172
rect 15929 14112 15993 14116
rect 16009 14172 16073 14176
rect 16009 14116 16013 14172
rect 16013 14116 16069 14172
rect 16069 14116 16073 14172
rect 16009 14112 16073 14116
rect 16089 14172 16153 14176
rect 16089 14116 16093 14172
rect 16093 14116 16149 14172
rect 16149 14116 16153 14172
rect 16089 14112 16153 14116
rect 16169 14172 16233 14176
rect 16169 14116 16173 14172
rect 16173 14116 16229 14172
rect 16229 14116 16233 14172
rect 16169 14112 16233 14116
rect 21656 14172 21720 14176
rect 21656 14116 21660 14172
rect 21660 14116 21716 14172
rect 21716 14116 21720 14172
rect 21656 14112 21720 14116
rect 21736 14172 21800 14176
rect 21736 14116 21740 14172
rect 21740 14116 21796 14172
rect 21796 14116 21800 14172
rect 21736 14112 21800 14116
rect 21816 14172 21880 14176
rect 21816 14116 21820 14172
rect 21820 14116 21876 14172
rect 21876 14116 21880 14172
rect 21816 14112 21880 14116
rect 21896 14172 21960 14176
rect 21896 14116 21900 14172
rect 21900 14116 21956 14172
rect 21956 14116 21960 14172
rect 21896 14112 21960 14116
rect 3815 13628 3879 13632
rect 3815 13572 3819 13628
rect 3819 13572 3875 13628
rect 3875 13572 3879 13628
rect 3815 13568 3879 13572
rect 3895 13628 3959 13632
rect 3895 13572 3899 13628
rect 3899 13572 3955 13628
rect 3955 13572 3959 13628
rect 3895 13568 3959 13572
rect 3975 13628 4039 13632
rect 3975 13572 3979 13628
rect 3979 13572 4035 13628
rect 4035 13572 4039 13628
rect 3975 13568 4039 13572
rect 4055 13628 4119 13632
rect 4055 13572 4059 13628
rect 4059 13572 4115 13628
rect 4115 13572 4119 13628
rect 4055 13568 4119 13572
rect 9542 13628 9606 13632
rect 9542 13572 9546 13628
rect 9546 13572 9602 13628
rect 9602 13572 9606 13628
rect 9542 13568 9606 13572
rect 9622 13628 9686 13632
rect 9622 13572 9626 13628
rect 9626 13572 9682 13628
rect 9682 13572 9686 13628
rect 9622 13568 9686 13572
rect 9702 13628 9766 13632
rect 9702 13572 9706 13628
rect 9706 13572 9762 13628
rect 9762 13572 9766 13628
rect 9702 13568 9766 13572
rect 9782 13628 9846 13632
rect 9782 13572 9786 13628
rect 9786 13572 9842 13628
rect 9842 13572 9846 13628
rect 9782 13568 9846 13572
rect 15269 13628 15333 13632
rect 15269 13572 15273 13628
rect 15273 13572 15329 13628
rect 15329 13572 15333 13628
rect 15269 13568 15333 13572
rect 15349 13628 15413 13632
rect 15349 13572 15353 13628
rect 15353 13572 15409 13628
rect 15409 13572 15413 13628
rect 15349 13568 15413 13572
rect 15429 13628 15493 13632
rect 15429 13572 15433 13628
rect 15433 13572 15489 13628
rect 15489 13572 15493 13628
rect 15429 13568 15493 13572
rect 15509 13628 15573 13632
rect 15509 13572 15513 13628
rect 15513 13572 15569 13628
rect 15569 13572 15573 13628
rect 15509 13568 15573 13572
rect 20996 13628 21060 13632
rect 20996 13572 21000 13628
rect 21000 13572 21056 13628
rect 21056 13572 21060 13628
rect 20996 13568 21060 13572
rect 21076 13628 21140 13632
rect 21076 13572 21080 13628
rect 21080 13572 21136 13628
rect 21136 13572 21140 13628
rect 21076 13568 21140 13572
rect 21156 13628 21220 13632
rect 21156 13572 21160 13628
rect 21160 13572 21216 13628
rect 21216 13572 21220 13628
rect 21156 13568 21220 13572
rect 21236 13628 21300 13632
rect 21236 13572 21240 13628
rect 21240 13572 21296 13628
rect 21296 13572 21300 13628
rect 21236 13568 21300 13572
rect 4475 13084 4539 13088
rect 4475 13028 4479 13084
rect 4479 13028 4535 13084
rect 4535 13028 4539 13084
rect 4475 13024 4539 13028
rect 4555 13084 4619 13088
rect 4555 13028 4559 13084
rect 4559 13028 4615 13084
rect 4615 13028 4619 13084
rect 4555 13024 4619 13028
rect 4635 13084 4699 13088
rect 4635 13028 4639 13084
rect 4639 13028 4695 13084
rect 4695 13028 4699 13084
rect 4635 13024 4699 13028
rect 4715 13084 4779 13088
rect 4715 13028 4719 13084
rect 4719 13028 4775 13084
rect 4775 13028 4779 13084
rect 4715 13024 4779 13028
rect 10202 13084 10266 13088
rect 10202 13028 10206 13084
rect 10206 13028 10262 13084
rect 10262 13028 10266 13084
rect 10202 13024 10266 13028
rect 10282 13084 10346 13088
rect 10282 13028 10286 13084
rect 10286 13028 10342 13084
rect 10342 13028 10346 13084
rect 10282 13024 10346 13028
rect 10362 13084 10426 13088
rect 10362 13028 10366 13084
rect 10366 13028 10422 13084
rect 10422 13028 10426 13084
rect 10362 13024 10426 13028
rect 10442 13084 10506 13088
rect 10442 13028 10446 13084
rect 10446 13028 10502 13084
rect 10502 13028 10506 13084
rect 10442 13024 10506 13028
rect 15929 13084 15993 13088
rect 15929 13028 15933 13084
rect 15933 13028 15989 13084
rect 15989 13028 15993 13084
rect 15929 13024 15993 13028
rect 16009 13084 16073 13088
rect 16009 13028 16013 13084
rect 16013 13028 16069 13084
rect 16069 13028 16073 13084
rect 16009 13024 16073 13028
rect 16089 13084 16153 13088
rect 16089 13028 16093 13084
rect 16093 13028 16149 13084
rect 16149 13028 16153 13084
rect 16089 13024 16153 13028
rect 16169 13084 16233 13088
rect 16169 13028 16173 13084
rect 16173 13028 16229 13084
rect 16229 13028 16233 13084
rect 16169 13024 16233 13028
rect 21656 13084 21720 13088
rect 21656 13028 21660 13084
rect 21660 13028 21716 13084
rect 21716 13028 21720 13084
rect 21656 13024 21720 13028
rect 21736 13084 21800 13088
rect 21736 13028 21740 13084
rect 21740 13028 21796 13084
rect 21796 13028 21800 13084
rect 21736 13024 21800 13028
rect 21816 13084 21880 13088
rect 21816 13028 21820 13084
rect 21820 13028 21876 13084
rect 21876 13028 21880 13084
rect 21816 13024 21880 13028
rect 21896 13084 21960 13088
rect 21896 13028 21900 13084
rect 21900 13028 21956 13084
rect 21956 13028 21960 13084
rect 21896 13024 21960 13028
rect 3815 12540 3879 12544
rect 3815 12484 3819 12540
rect 3819 12484 3875 12540
rect 3875 12484 3879 12540
rect 3815 12480 3879 12484
rect 3895 12540 3959 12544
rect 3895 12484 3899 12540
rect 3899 12484 3955 12540
rect 3955 12484 3959 12540
rect 3895 12480 3959 12484
rect 3975 12540 4039 12544
rect 3975 12484 3979 12540
rect 3979 12484 4035 12540
rect 4035 12484 4039 12540
rect 3975 12480 4039 12484
rect 4055 12540 4119 12544
rect 4055 12484 4059 12540
rect 4059 12484 4115 12540
rect 4115 12484 4119 12540
rect 4055 12480 4119 12484
rect 9542 12540 9606 12544
rect 9542 12484 9546 12540
rect 9546 12484 9602 12540
rect 9602 12484 9606 12540
rect 9542 12480 9606 12484
rect 9622 12540 9686 12544
rect 9622 12484 9626 12540
rect 9626 12484 9682 12540
rect 9682 12484 9686 12540
rect 9622 12480 9686 12484
rect 9702 12540 9766 12544
rect 9702 12484 9706 12540
rect 9706 12484 9762 12540
rect 9762 12484 9766 12540
rect 9702 12480 9766 12484
rect 9782 12540 9846 12544
rect 9782 12484 9786 12540
rect 9786 12484 9842 12540
rect 9842 12484 9846 12540
rect 9782 12480 9846 12484
rect 15269 12540 15333 12544
rect 15269 12484 15273 12540
rect 15273 12484 15329 12540
rect 15329 12484 15333 12540
rect 15269 12480 15333 12484
rect 15349 12540 15413 12544
rect 15349 12484 15353 12540
rect 15353 12484 15409 12540
rect 15409 12484 15413 12540
rect 15349 12480 15413 12484
rect 15429 12540 15493 12544
rect 15429 12484 15433 12540
rect 15433 12484 15489 12540
rect 15489 12484 15493 12540
rect 15429 12480 15493 12484
rect 15509 12540 15573 12544
rect 15509 12484 15513 12540
rect 15513 12484 15569 12540
rect 15569 12484 15573 12540
rect 15509 12480 15573 12484
rect 20996 12540 21060 12544
rect 20996 12484 21000 12540
rect 21000 12484 21056 12540
rect 21056 12484 21060 12540
rect 20996 12480 21060 12484
rect 21076 12540 21140 12544
rect 21076 12484 21080 12540
rect 21080 12484 21136 12540
rect 21136 12484 21140 12540
rect 21076 12480 21140 12484
rect 21156 12540 21220 12544
rect 21156 12484 21160 12540
rect 21160 12484 21216 12540
rect 21216 12484 21220 12540
rect 21156 12480 21220 12484
rect 21236 12540 21300 12544
rect 21236 12484 21240 12540
rect 21240 12484 21296 12540
rect 21296 12484 21300 12540
rect 21236 12480 21300 12484
rect 4475 11996 4539 12000
rect 4475 11940 4479 11996
rect 4479 11940 4535 11996
rect 4535 11940 4539 11996
rect 4475 11936 4539 11940
rect 4555 11996 4619 12000
rect 4555 11940 4559 11996
rect 4559 11940 4615 11996
rect 4615 11940 4619 11996
rect 4555 11936 4619 11940
rect 4635 11996 4699 12000
rect 4635 11940 4639 11996
rect 4639 11940 4695 11996
rect 4695 11940 4699 11996
rect 4635 11936 4699 11940
rect 4715 11996 4779 12000
rect 4715 11940 4719 11996
rect 4719 11940 4775 11996
rect 4775 11940 4779 11996
rect 4715 11936 4779 11940
rect 10202 11996 10266 12000
rect 10202 11940 10206 11996
rect 10206 11940 10262 11996
rect 10262 11940 10266 11996
rect 10202 11936 10266 11940
rect 10282 11996 10346 12000
rect 10282 11940 10286 11996
rect 10286 11940 10342 11996
rect 10342 11940 10346 11996
rect 10282 11936 10346 11940
rect 10362 11996 10426 12000
rect 10362 11940 10366 11996
rect 10366 11940 10422 11996
rect 10422 11940 10426 11996
rect 10362 11936 10426 11940
rect 10442 11996 10506 12000
rect 10442 11940 10446 11996
rect 10446 11940 10502 11996
rect 10502 11940 10506 11996
rect 10442 11936 10506 11940
rect 15929 11996 15993 12000
rect 15929 11940 15933 11996
rect 15933 11940 15989 11996
rect 15989 11940 15993 11996
rect 15929 11936 15993 11940
rect 16009 11996 16073 12000
rect 16009 11940 16013 11996
rect 16013 11940 16069 11996
rect 16069 11940 16073 11996
rect 16009 11936 16073 11940
rect 16089 11996 16153 12000
rect 16089 11940 16093 11996
rect 16093 11940 16149 11996
rect 16149 11940 16153 11996
rect 16089 11936 16153 11940
rect 16169 11996 16233 12000
rect 16169 11940 16173 11996
rect 16173 11940 16229 11996
rect 16229 11940 16233 11996
rect 16169 11936 16233 11940
rect 21656 11996 21720 12000
rect 21656 11940 21660 11996
rect 21660 11940 21716 11996
rect 21716 11940 21720 11996
rect 21656 11936 21720 11940
rect 21736 11996 21800 12000
rect 21736 11940 21740 11996
rect 21740 11940 21796 11996
rect 21796 11940 21800 11996
rect 21736 11936 21800 11940
rect 21816 11996 21880 12000
rect 21816 11940 21820 11996
rect 21820 11940 21876 11996
rect 21876 11940 21880 11996
rect 21816 11936 21880 11940
rect 21896 11996 21960 12000
rect 21896 11940 21900 11996
rect 21900 11940 21956 11996
rect 21956 11940 21960 11996
rect 21896 11936 21960 11940
rect 3815 11452 3879 11456
rect 3815 11396 3819 11452
rect 3819 11396 3875 11452
rect 3875 11396 3879 11452
rect 3815 11392 3879 11396
rect 3895 11452 3959 11456
rect 3895 11396 3899 11452
rect 3899 11396 3955 11452
rect 3955 11396 3959 11452
rect 3895 11392 3959 11396
rect 3975 11452 4039 11456
rect 3975 11396 3979 11452
rect 3979 11396 4035 11452
rect 4035 11396 4039 11452
rect 3975 11392 4039 11396
rect 4055 11452 4119 11456
rect 4055 11396 4059 11452
rect 4059 11396 4115 11452
rect 4115 11396 4119 11452
rect 4055 11392 4119 11396
rect 9542 11452 9606 11456
rect 9542 11396 9546 11452
rect 9546 11396 9602 11452
rect 9602 11396 9606 11452
rect 9542 11392 9606 11396
rect 9622 11452 9686 11456
rect 9622 11396 9626 11452
rect 9626 11396 9682 11452
rect 9682 11396 9686 11452
rect 9622 11392 9686 11396
rect 9702 11452 9766 11456
rect 9702 11396 9706 11452
rect 9706 11396 9762 11452
rect 9762 11396 9766 11452
rect 9702 11392 9766 11396
rect 9782 11452 9846 11456
rect 9782 11396 9786 11452
rect 9786 11396 9842 11452
rect 9842 11396 9846 11452
rect 9782 11392 9846 11396
rect 15269 11452 15333 11456
rect 15269 11396 15273 11452
rect 15273 11396 15329 11452
rect 15329 11396 15333 11452
rect 15269 11392 15333 11396
rect 15349 11452 15413 11456
rect 15349 11396 15353 11452
rect 15353 11396 15409 11452
rect 15409 11396 15413 11452
rect 15349 11392 15413 11396
rect 15429 11452 15493 11456
rect 15429 11396 15433 11452
rect 15433 11396 15489 11452
rect 15489 11396 15493 11452
rect 15429 11392 15493 11396
rect 15509 11452 15573 11456
rect 15509 11396 15513 11452
rect 15513 11396 15569 11452
rect 15569 11396 15573 11452
rect 15509 11392 15573 11396
rect 20996 11452 21060 11456
rect 20996 11396 21000 11452
rect 21000 11396 21056 11452
rect 21056 11396 21060 11452
rect 20996 11392 21060 11396
rect 21076 11452 21140 11456
rect 21076 11396 21080 11452
rect 21080 11396 21136 11452
rect 21136 11396 21140 11452
rect 21076 11392 21140 11396
rect 21156 11452 21220 11456
rect 21156 11396 21160 11452
rect 21160 11396 21216 11452
rect 21216 11396 21220 11452
rect 21156 11392 21220 11396
rect 21236 11452 21300 11456
rect 21236 11396 21240 11452
rect 21240 11396 21296 11452
rect 21296 11396 21300 11452
rect 21236 11392 21300 11396
rect 4475 10908 4539 10912
rect 4475 10852 4479 10908
rect 4479 10852 4535 10908
rect 4535 10852 4539 10908
rect 4475 10848 4539 10852
rect 4555 10908 4619 10912
rect 4555 10852 4559 10908
rect 4559 10852 4615 10908
rect 4615 10852 4619 10908
rect 4555 10848 4619 10852
rect 4635 10908 4699 10912
rect 4635 10852 4639 10908
rect 4639 10852 4695 10908
rect 4695 10852 4699 10908
rect 4635 10848 4699 10852
rect 4715 10908 4779 10912
rect 4715 10852 4719 10908
rect 4719 10852 4775 10908
rect 4775 10852 4779 10908
rect 4715 10848 4779 10852
rect 10202 10908 10266 10912
rect 10202 10852 10206 10908
rect 10206 10852 10262 10908
rect 10262 10852 10266 10908
rect 10202 10848 10266 10852
rect 10282 10908 10346 10912
rect 10282 10852 10286 10908
rect 10286 10852 10342 10908
rect 10342 10852 10346 10908
rect 10282 10848 10346 10852
rect 10362 10908 10426 10912
rect 10362 10852 10366 10908
rect 10366 10852 10422 10908
rect 10422 10852 10426 10908
rect 10362 10848 10426 10852
rect 10442 10908 10506 10912
rect 10442 10852 10446 10908
rect 10446 10852 10502 10908
rect 10502 10852 10506 10908
rect 10442 10848 10506 10852
rect 15929 10908 15993 10912
rect 15929 10852 15933 10908
rect 15933 10852 15989 10908
rect 15989 10852 15993 10908
rect 15929 10848 15993 10852
rect 16009 10908 16073 10912
rect 16009 10852 16013 10908
rect 16013 10852 16069 10908
rect 16069 10852 16073 10908
rect 16009 10848 16073 10852
rect 16089 10908 16153 10912
rect 16089 10852 16093 10908
rect 16093 10852 16149 10908
rect 16149 10852 16153 10908
rect 16089 10848 16153 10852
rect 16169 10908 16233 10912
rect 16169 10852 16173 10908
rect 16173 10852 16229 10908
rect 16229 10852 16233 10908
rect 16169 10848 16233 10852
rect 21656 10908 21720 10912
rect 21656 10852 21660 10908
rect 21660 10852 21716 10908
rect 21716 10852 21720 10908
rect 21656 10848 21720 10852
rect 21736 10908 21800 10912
rect 21736 10852 21740 10908
rect 21740 10852 21796 10908
rect 21796 10852 21800 10908
rect 21736 10848 21800 10852
rect 21816 10908 21880 10912
rect 21816 10852 21820 10908
rect 21820 10852 21876 10908
rect 21876 10852 21880 10908
rect 21816 10848 21880 10852
rect 21896 10908 21960 10912
rect 21896 10852 21900 10908
rect 21900 10852 21956 10908
rect 21956 10852 21960 10908
rect 21896 10848 21960 10852
rect 3815 10364 3879 10368
rect 3815 10308 3819 10364
rect 3819 10308 3875 10364
rect 3875 10308 3879 10364
rect 3815 10304 3879 10308
rect 3895 10364 3959 10368
rect 3895 10308 3899 10364
rect 3899 10308 3955 10364
rect 3955 10308 3959 10364
rect 3895 10304 3959 10308
rect 3975 10364 4039 10368
rect 3975 10308 3979 10364
rect 3979 10308 4035 10364
rect 4035 10308 4039 10364
rect 3975 10304 4039 10308
rect 4055 10364 4119 10368
rect 4055 10308 4059 10364
rect 4059 10308 4115 10364
rect 4115 10308 4119 10364
rect 4055 10304 4119 10308
rect 9542 10364 9606 10368
rect 9542 10308 9546 10364
rect 9546 10308 9602 10364
rect 9602 10308 9606 10364
rect 9542 10304 9606 10308
rect 9622 10364 9686 10368
rect 9622 10308 9626 10364
rect 9626 10308 9682 10364
rect 9682 10308 9686 10364
rect 9622 10304 9686 10308
rect 9702 10364 9766 10368
rect 9702 10308 9706 10364
rect 9706 10308 9762 10364
rect 9762 10308 9766 10364
rect 9702 10304 9766 10308
rect 9782 10364 9846 10368
rect 9782 10308 9786 10364
rect 9786 10308 9842 10364
rect 9842 10308 9846 10364
rect 9782 10304 9846 10308
rect 15269 10364 15333 10368
rect 15269 10308 15273 10364
rect 15273 10308 15329 10364
rect 15329 10308 15333 10364
rect 15269 10304 15333 10308
rect 15349 10364 15413 10368
rect 15349 10308 15353 10364
rect 15353 10308 15409 10364
rect 15409 10308 15413 10364
rect 15349 10304 15413 10308
rect 15429 10364 15493 10368
rect 15429 10308 15433 10364
rect 15433 10308 15489 10364
rect 15489 10308 15493 10364
rect 15429 10304 15493 10308
rect 15509 10364 15573 10368
rect 15509 10308 15513 10364
rect 15513 10308 15569 10364
rect 15569 10308 15573 10364
rect 15509 10304 15573 10308
rect 20996 10364 21060 10368
rect 20996 10308 21000 10364
rect 21000 10308 21056 10364
rect 21056 10308 21060 10364
rect 20996 10304 21060 10308
rect 21076 10364 21140 10368
rect 21076 10308 21080 10364
rect 21080 10308 21136 10364
rect 21136 10308 21140 10364
rect 21076 10304 21140 10308
rect 21156 10364 21220 10368
rect 21156 10308 21160 10364
rect 21160 10308 21216 10364
rect 21216 10308 21220 10364
rect 21156 10304 21220 10308
rect 21236 10364 21300 10368
rect 21236 10308 21240 10364
rect 21240 10308 21296 10364
rect 21296 10308 21300 10364
rect 21236 10304 21300 10308
rect 4475 9820 4539 9824
rect 4475 9764 4479 9820
rect 4479 9764 4535 9820
rect 4535 9764 4539 9820
rect 4475 9760 4539 9764
rect 4555 9820 4619 9824
rect 4555 9764 4559 9820
rect 4559 9764 4615 9820
rect 4615 9764 4619 9820
rect 4555 9760 4619 9764
rect 4635 9820 4699 9824
rect 4635 9764 4639 9820
rect 4639 9764 4695 9820
rect 4695 9764 4699 9820
rect 4635 9760 4699 9764
rect 4715 9820 4779 9824
rect 4715 9764 4719 9820
rect 4719 9764 4775 9820
rect 4775 9764 4779 9820
rect 4715 9760 4779 9764
rect 10202 9820 10266 9824
rect 10202 9764 10206 9820
rect 10206 9764 10262 9820
rect 10262 9764 10266 9820
rect 10202 9760 10266 9764
rect 10282 9820 10346 9824
rect 10282 9764 10286 9820
rect 10286 9764 10342 9820
rect 10342 9764 10346 9820
rect 10282 9760 10346 9764
rect 10362 9820 10426 9824
rect 10362 9764 10366 9820
rect 10366 9764 10422 9820
rect 10422 9764 10426 9820
rect 10362 9760 10426 9764
rect 10442 9820 10506 9824
rect 10442 9764 10446 9820
rect 10446 9764 10502 9820
rect 10502 9764 10506 9820
rect 10442 9760 10506 9764
rect 15929 9820 15993 9824
rect 15929 9764 15933 9820
rect 15933 9764 15989 9820
rect 15989 9764 15993 9820
rect 15929 9760 15993 9764
rect 16009 9820 16073 9824
rect 16009 9764 16013 9820
rect 16013 9764 16069 9820
rect 16069 9764 16073 9820
rect 16009 9760 16073 9764
rect 16089 9820 16153 9824
rect 16089 9764 16093 9820
rect 16093 9764 16149 9820
rect 16149 9764 16153 9820
rect 16089 9760 16153 9764
rect 16169 9820 16233 9824
rect 16169 9764 16173 9820
rect 16173 9764 16229 9820
rect 16229 9764 16233 9820
rect 16169 9760 16233 9764
rect 21656 9820 21720 9824
rect 21656 9764 21660 9820
rect 21660 9764 21716 9820
rect 21716 9764 21720 9820
rect 21656 9760 21720 9764
rect 21736 9820 21800 9824
rect 21736 9764 21740 9820
rect 21740 9764 21796 9820
rect 21796 9764 21800 9820
rect 21736 9760 21800 9764
rect 21816 9820 21880 9824
rect 21816 9764 21820 9820
rect 21820 9764 21876 9820
rect 21876 9764 21880 9820
rect 21816 9760 21880 9764
rect 21896 9820 21960 9824
rect 21896 9764 21900 9820
rect 21900 9764 21956 9820
rect 21956 9764 21960 9820
rect 21896 9760 21960 9764
rect 3815 9276 3879 9280
rect 3815 9220 3819 9276
rect 3819 9220 3875 9276
rect 3875 9220 3879 9276
rect 3815 9216 3879 9220
rect 3895 9276 3959 9280
rect 3895 9220 3899 9276
rect 3899 9220 3955 9276
rect 3955 9220 3959 9276
rect 3895 9216 3959 9220
rect 3975 9276 4039 9280
rect 3975 9220 3979 9276
rect 3979 9220 4035 9276
rect 4035 9220 4039 9276
rect 3975 9216 4039 9220
rect 4055 9276 4119 9280
rect 4055 9220 4059 9276
rect 4059 9220 4115 9276
rect 4115 9220 4119 9276
rect 4055 9216 4119 9220
rect 9542 9276 9606 9280
rect 9542 9220 9546 9276
rect 9546 9220 9602 9276
rect 9602 9220 9606 9276
rect 9542 9216 9606 9220
rect 9622 9276 9686 9280
rect 9622 9220 9626 9276
rect 9626 9220 9682 9276
rect 9682 9220 9686 9276
rect 9622 9216 9686 9220
rect 9702 9276 9766 9280
rect 9702 9220 9706 9276
rect 9706 9220 9762 9276
rect 9762 9220 9766 9276
rect 9702 9216 9766 9220
rect 9782 9276 9846 9280
rect 9782 9220 9786 9276
rect 9786 9220 9842 9276
rect 9842 9220 9846 9276
rect 9782 9216 9846 9220
rect 15269 9276 15333 9280
rect 15269 9220 15273 9276
rect 15273 9220 15329 9276
rect 15329 9220 15333 9276
rect 15269 9216 15333 9220
rect 15349 9276 15413 9280
rect 15349 9220 15353 9276
rect 15353 9220 15409 9276
rect 15409 9220 15413 9276
rect 15349 9216 15413 9220
rect 15429 9276 15493 9280
rect 15429 9220 15433 9276
rect 15433 9220 15489 9276
rect 15489 9220 15493 9276
rect 15429 9216 15493 9220
rect 15509 9276 15573 9280
rect 15509 9220 15513 9276
rect 15513 9220 15569 9276
rect 15569 9220 15573 9276
rect 15509 9216 15573 9220
rect 20996 9276 21060 9280
rect 20996 9220 21000 9276
rect 21000 9220 21056 9276
rect 21056 9220 21060 9276
rect 20996 9216 21060 9220
rect 21076 9276 21140 9280
rect 21076 9220 21080 9276
rect 21080 9220 21136 9276
rect 21136 9220 21140 9276
rect 21076 9216 21140 9220
rect 21156 9276 21220 9280
rect 21156 9220 21160 9276
rect 21160 9220 21216 9276
rect 21216 9220 21220 9276
rect 21156 9216 21220 9220
rect 21236 9276 21300 9280
rect 21236 9220 21240 9276
rect 21240 9220 21296 9276
rect 21296 9220 21300 9276
rect 21236 9216 21300 9220
rect 4475 8732 4539 8736
rect 4475 8676 4479 8732
rect 4479 8676 4535 8732
rect 4535 8676 4539 8732
rect 4475 8672 4539 8676
rect 4555 8732 4619 8736
rect 4555 8676 4559 8732
rect 4559 8676 4615 8732
rect 4615 8676 4619 8732
rect 4555 8672 4619 8676
rect 4635 8732 4699 8736
rect 4635 8676 4639 8732
rect 4639 8676 4695 8732
rect 4695 8676 4699 8732
rect 4635 8672 4699 8676
rect 4715 8732 4779 8736
rect 4715 8676 4719 8732
rect 4719 8676 4775 8732
rect 4775 8676 4779 8732
rect 4715 8672 4779 8676
rect 10202 8732 10266 8736
rect 10202 8676 10206 8732
rect 10206 8676 10262 8732
rect 10262 8676 10266 8732
rect 10202 8672 10266 8676
rect 10282 8732 10346 8736
rect 10282 8676 10286 8732
rect 10286 8676 10342 8732
rect 10342 8676 10346 8732
rect 10282 8672 10346 8676
rect 10362 8732 10426 8736
rect 10362 8676 10366 8732
rect 10366 8676 10422 8732
rect 10422 8676 10426 8732
rect 10362 8672 10426 8676
rect 10442 8732 10506 8736
rect 10442 8676 10446 8732
rect 10446 8676 10502 8732
rect 10502 8676 10506 8732
rect 10442 8672 10506 8676
rect 15929 8732 15993 8736
rect 15929 8676 15933 8732
rect 15933 8676 15989 8732
rect 15989 8676 15993 8732
rect 15929 8672 15993 8676
rect 16009 8732 16073 8736
rect 16009 8676 16013 8732
rect 16013 8676 16069 8732
rect 16069 8676 16073 8732
rect 16009 8672 16073 8676
rect 16089 8732 16153 8736
rect 16089 8676 16093 8732
rect 16093 8676 16149 8732
rect 16149 8676 16153 8732
rect 16089 8672 16153 8676
rect 16169 8732 16233 8736
rect 16169 8676 16173 8732
rect 16173 8676 16229 8732
rect 16229 8676 16233 8732
rect 16169 8672 16233 8676
rect 21656 8732 21720 8736
rect 21656 8676 21660 8732
rect 21660 8676 21716 8732
rect 21716 8676 21720 8732
rect 21656 8672 21720 8676
rect 21736 8732 21800 8736
rect 21736 8676 21740 8732
rect 21740 8676 21796 8732
rect 21796 8676 21800 8732
rect 21736 8672 21800 8676
rect 21816 8732 21880 8736
rect 21816 8676 21820 8732
rect 21820 8676 21876 8732
rect 21876 8676 21880 8732
rect 21816 8672 21880 8676
rect 21896 8732 21960 8736
rect 21896 8676 21900 8732
rect 21900 8676 21956 8732
rect 21956 8676 21960 8732
rect 21896 8672 21960 8676
rect 3815 8188 3879 8192
rect 3815 8132 3819 8188
rect 3819 8132 3875 8188
rect 3875 8132 3879 8188
rect 3815 8128 3879 8132
rect 3895 8188 3959 8192
rect 3895 8132 3899 8188
rect 3899 8132 3955 8188
rect 3955 8132 3959 8188
rect 3895 8128 3959 8132
rect 3975 8188 4039 8192
rect 3975 8132 3979 8188
rect 3979 8132 4035 8188
rect 4035 8132 4039 8188
rect 3975 8128 4039 8132
rect 4055 8188 4119 8192
rect 4055 8132 4059 8188
rect 4059 8132 4115 8188
rect 4115 8132 4119 8188
rect 4055 8128 4119 8132
rect 9542 8188 9606 8192
rect 9542 8132 9546 8188
rect 9546 8132 9602 8188
rect 9602 8132 9606 8188
rect 9542 8128 9606 8132
rect 9622 8188 9686 8192
rect 9622 8132 9626 8188
rect 9626 8132 9682 8188
rect 9682 8132 9686 8188
rect 9622 8128 9686 8132
rect 9702 8188 9766 8192
rect 9702 8132 9706 8188
rect 9706 8132 9762 8188
rect 9762 8132 9766 8188
rect 9702 8128 9766 8132
rect 9782 8188 9846 8192
rect 9782 8132 9786 8188
rect 9786 8132 9842 8188
rect 9842 8132 9846 8188
rect 9782 8128 9846 8132
rect 15269 8188 15333 8192
rect 15269 8132 15273 8188
rect 15273 8132 15329 8188
rect 15329 8132 15333 8188
rect 15269 8128 15333 8132
rect 15349 8188 15413 8192
rect 15349 8132 15353 8188
rect 15353 8132 15409 8188
rect 15409 8132 15413 8188
rect 15349 8128 15413 8132
rect 15429 8188 15493 8192
rect 15429 8132 15433 8188
rect 15433 8132 15489 8188
rect 15489 8132 15493 8188
rect 15429 8128 15493 8132
rect 15509 8188 15573 8192
rect 15509 8132 15513 8188
rect 15513 8132 15569 8188
rect 15569 8132 15573 8188
rect 15509 8128 15573 8132
rect 20996 8188 21060 8192
rect 20996 8132 21000 8188
rect 21000 8132 21056 8188
rect 21056 8132 21060 8188
rect 20996 8128 21060 8132
rect 21076 8188 21140 8192
rect 21076 8132 21080 8188
rect 21080 8132 21136 8188
rect 21136 8132 21140 8188
rect 21076 8128 21140 8132
rect 21156 8188 21220 8192
rect 21156 8132 21160 8188
rect 21160 8132 21216 8188
rect 21216 8132 21220 8188
rect 21156 8128 21220 8132
rect 21236 8188 21300 8192
rect 21236 8132 21240 8188
rect 21240 8132 21296 8188
rect 21296 8132 21300 8188
rect 21236 8128 21300 8132
rect 4475 7644 4539 7648
rect 4475 7588 4479 7644
rect 4479 7588 4535 7644
rect 4535 7588 4539 7644
rect 4475 7584 4539 7588
rect 4555 7644 4619 7648
rect 4555 7588 4559 7644
rect 4559 7588 4615 7644
rect 4615 7588 4619 7644
rect 4555 7584 4619 7588
rect 4635 7644 4699 7648
rect 4635 7588 4639 7644
rect 4639 7588 4695 7644
rect 4695 7588 4699 7644
rect 4635 7584 4699 7588
rect 4715 7644 4779 7648
rect 4715 7588 4719 7644
rect 4719 7588 4775 7644
rect 4775 7588 4779 7644
rect 4715 7584 4779 7588
rect 10202 7644 10266 7648
rect 10202 7588 10206 7644
rect 10206 7588 10262 7644
rect 10262 7588 10266 7644
rect 10202 7584 10266 7588
rect 10282 7644 10346 7648
rect 10282 7588 10286 7644
rect 10286 7588 10342 7644
rect 10342 7588 10346 7644
rect 10282 7584 10346 7588
rect 10362 7644 10426 7648
rect 10362 7588 10366 7644
rect 10366 7588 10422 7644
rect 10422 7588 10426 7644
rect 10362 7584 10426 7588
rect 10442 7644 10506 7648
rect 10442 7588 10446 7644
rect 10446 7588 10502 7644
rect 10502 7588 10506 7644
rect 10442 7584 10506 7588
rect 15929 7644 15993 7648
rect 15929 7588 15933 7644
rect 15933 7588 15989 7644
rect 15989 7588 15993 7644
rect 15929 7584 15993 7588
rect 16009 7644 16073 7648
rect 16009 7588 16013 7644
rect 16013 7588 16069 7644
rect 16069 7588 16073 7644
rect 16009 7584 16073 7588
rect 16089 7644 16153 7648
rect 16089 7588 16093 7644
rect 16093 7588 16149 7644
rect 16149 7588 16153 7644
rect 16089 7584 16153 7588
rect 16169 7644 16233 7648
rect 16169 7588 16173 7644
rect 16173 7588 16229 7644
rect 16229 7588 16233 7644
rect 16169 7584 16233 7588
rect 21656 7644 21720 7648
rect 21656 7588 21660 7644
rect 21660 7588 21716 7644
rect 21716 7588 21720 7644
rect 21656 7584 21720 7588
rect 21736 7644 21800 7648
rect 21736 7588 21740 7644
rect 21740 7588 21796 7644
rect 21796 7588 21800 7644
rect 21736 7584 21800 7588
rect 21816 7644 21880 7648
rect 21816 7588 21820 7644
rect 21820 7588 21876 7644
rect 21876 7588 21880 7644
rect 21816 7584 21880 7588
rect 21896 7644 21960 7648
rect 21896 7588 21900 7644
rect 21900 7588 21956 7644
rect 21956 7588 21960 7644
rect 21896 7584 21960 7588
rect 3815 7100 3879 7104
rect 3815 7044 3819 7100
rect 3819 7044 3875 7100
rect 3875 7044 3879 7100
rect 3815 7040 3879 7044
rect 3895 7100 3959 7104
rect 3895 7044 3899 7100
rect 3899 7044 3955 7100
rect 3955 7044 3959 7100
rect 3895 7040 3959 7044
rect 3975 7100 4039 7104
rect 3975 7044 3979 7100
rect 3979 7044 4035 7100
rect 4035 7044 4039 7100
rect 3975 7040 4039 7044
rect 4055 7100 4119 7104
rect 4055 7044 4059 7100
rect 4059 7044 4115 7100
rect 4115 7044 4119 7100
rect 4055 7040 4119 7044
rect 9542 7100 9606 7104
rect 9542 7044 9546 7100
rect 9546 7044 9602 7100
rect 9602 7044 9606 7100
rect 9542 7040 9606 7044
rect 9622 7100 9686 7104
rect 9622 7044 9626 7100
rect 9626 7044 9682 7100
rect 9682 7044 9686 7100
rect 9622 7040 9686 7044
rect 9702 7100 9766 7104
rect 9702 7044 9706 7100
rect 9706 7044 9762 7100
rect 9762 7044 9766 7100
rect 9702 7040 9766 7044
rect 9782 7100 9846 7104
rect 9782 7044 9786 7100
rect 9786 7044 9842 7100
rect 9842 7044 9846 7100
rect 9782 7040 9846 7044
rect 15269 7100 15333 7104
rect 15269 7044 15273 7100
rect 15273 7044 15329 7100
rect 15329 7044 15333 7100
rect 15269 7040 15333 7044
rect 15349 7100 15413 7104
rect 15349 7044 15353 7100
rect 15353 7044 15409 7100
rect 15409 7044 15413 7100
rect 15349 7040 15413 7044
rect 15429 7100 15493 7104
rect 15429 7044 15433 7100
rect 15433 7044 15489 7100
rect 15489 7044 15493 7100
rect 15429 7040 15493 7044
rect 15509 7100 15573 7104
rect 15509 7044 15513 7100
rect 15513 7044 15569 7100
rect 15569 7044 15573 7100
rect 15509 7040 15573 7044
rect 20996 7100 21060 7104
rect 20996 7044 21000 7100
rect 21000 7044 21056 7100
rect 21056 7044 21060 7100
rect 20996 7040 21060 7044
rect 21076 7100 21140 7104
rect 21076 7044 21080 7100
rect 21080 7044 21136 7100
rect 21136 7044 21140 7100
rect 21076 7040 21140 7044
rect 21156 7100 21220 7104
rect 21156 7044 21160 7100
rect 21160 7044 21216 7100
rect 21216 7044 21220 7100
rect 21156 7040 21220 7044
rect 21236 7100 21300 7104
rect 21236 7044 21240 7100
rect 21240 7044 21296 7100
rect 21296 7044 21300 7100
rect 21236 7040 21300 7044
rect 4475 6556 4539 6560
rect 4475 6500 4479 6556
rect 4479 6500 4535 6556
rect 4535 6500 4539 6556
rect 4475 6496 4539 6500
rect 4555 6556 4619 6560
rect 4555 6500 4559 6556
rect 4559 6500 4615 6556
rect 4615 6500 4619 6556
rect 4555 6496 4619 6500
rect 4635 6556 4699 6560
rect 4635 6500 4639 6556
rect 4639 6500 4695 6556
rect 4695 6500 4699 6556
rect 4635 6496 4699 6500
rect 4715 6556 4779 6560
rect 4715 6500 4719 6556
rect 4719 6500 4775 6556
rect 4775 6500 4779 6556
rect 4715 6496 4779 6500
rect 10202 6556 10266 6560
rect 10202 6500 10206 6556
rect 10206 6500 10262 6556
rect 10262 6500 10266 6556
rect 10202 6496 10266 6500
rect 10282 6556 10346 6560
rect 10282 6500 10286 6556
rect 10286 6500 10342 6556
rect 10342 6500 10346 6556
rect 10282 6496 10346 6500
rect 10362 6556 10426 6560
rect 10362 6500 10366 6556
rect 10366 6500 10422 6556
rect 10422 6500 10426 6556
rect 10362 6496 10426 6500
rect 10442 6556 10506 6560
rect 10442 6500 10446 6556
rect 10446 6500 10502 6556
rect 10502 6500 10506 6556
rect 10442 6496 10506 6500
rect 15929 6556 15993 6560
rect 15929 6500 15933 6556
rect 15933 6500 15989 6556
rect 15989 6500 15993 6556
rect 15929 6496 15993 6500
rect 16009 6556 16073 6560
rect 16009 6500 16013 6556
rect 16013 6500 16069 6556
rect 16069 6500 16073 6556
rect 16009 6496 16073 6500
rect 16089 6556 16153 6560
rect 16089 6500 16093 6556
rect 16093 6500 16149 6556
rect 16149 6500 16153 6556
rect 16089 6496 16153 6500
rect 16169 6556 16233 6560
rect 16169 6500 16173 6556
rect 16173 6500 16229 6556
rect 16229 6500 16233 6556
rect 16169 6496 16233 6500
rect 21656 6556 21720 6560
rect 21656 6500 21660 6556
rect 21660 6500 21716 6556
rect 21716 6500 21720 6556
rect 21656 6496 21720 6500
rect 21736 6556 21800 6560
rect 21736 6500 21740 6556
rect 21740 6500 21796 6556
rect 21796 6500 21800 6556
rect 21736 6496 21800 6500
rect 21816 6556 21880 6560
rect 21816 6500 21820 6556
rect 21820 6500 21876 6556
rect 21876 6500 21880 6556
rect 21816 6496 21880 6500
rect 21896 6556 21960 6560
rect 21896 6500 21900 6556
rect 21900 6500 21956 6556
rect 21956 6500 21960 6556
rect 21896 6496 21960 6500
rect 3815 6012 3879 6016
rect 3815 5956 3819 6012
rect 3819 5956 3875 6012
rect 3875 5956 3879 6012
rect 3815 5952 3879 5956
rect 3895 6012 3959 6016
rect 3895 5956 3899 6012
rect 3899 5956 3955 6012
rect 3955 5956 3959 6012
rect 3895 5952 3959 5956
rect 3975 6012 4039 6016
rect 3975 5956 3979 6012
rect 3979 5956 4035 6012
rect 4035 5956 4039 6012
rect 3975 5952 4039 5956
rect 4055 6012 4119 6016
rect 4055 5956 4059 6012
rect 4059 5956 4115 6012
rect 4115 5956 4119 6012
rect 4055 5952 4119 5956
rect 9542 6012 9606 6016
rect 9542 5956 9546 6012
rect 9546 5956 9602 6012
rect 9602 5956 9606 6012
rect 9542 5952 9606 5956
rect 9622 6012 9686 6016
rect 9622 5956 9626 6012
rect 9626 5956 9682 6012
rect 9682 5956 9686 6012
rect 9622 5952 9686 5956
rect 9702 6012 9766 6016
rect 9702 5956 9706 6012
rect 9706 5956 9762 6012
rect 9762 5956 9766 6012
rect 9702 5952 9766 5956
rect 9782 6012 9846 6016
rect 9782 5956 9786 6012
rect 9786 5956 9842 6012
rect 9842 5956 9846 6012
rect 9782 5952 9846 5956
rect 15269 6012 15333 6016
rect 15269 5956 15273 6012
rect 15273 5956 15329 6012
rect 15329 5956 15333 6012
rect 15269 5952 15333 5956
rect 15349 6012 15413 6016
rect 15349 5956 15353 6012
rect 15353 5956 15409 6012
rect 15409 5956 15413 6012
rect 15349 5952 15413 5956
rect 15429 6012 15493 6016
rect 15429 5956 15433 6012
rect 15433 5956 15489 6012
rect 15489 5956 15493 6012
rect 15429 5952 15493 5956
rect 15509 6012 15573 6016
rect 15509 5956 15513 6012
rect 15513 5956 15569 6012
rect 15569 5956 15573 6012
rect 15509 5952 15573 5956
rect 20996 6012 21060 6016
rect 20996 5956 21000 6012
rect 21000 5956 21056 6012
rect 21056 5956 21060 6012
rect 20996 5952 21060 5956
rect 21076 6012 21140 6016
rect 21076 5956 21080 6012
rect 21080 5956 21136 6012
rect 21136 5956 21140 6012
rect 21076 5952 21140 5956
rect 21156 6012 21220 6016
rect 21156 5956 21160 6012
rect 21160 5956 21216 6012
rect 21216 5956 21220 6012
rect 21156 5952 21220 5956
rect 21236 6012 21300 6016
rect 21236 5956 21240 6012
rect 21240 5956 21296 6012
rect 21296 5956 21300 6012
rect 21236 5952 21300 5956
rect 4475 5468 4539 5472
rect 4475 5412 4479 5468
rect 4479 5412 4535 5468
rect 4535 5412 4539 5468
rect 4475 5408 4539 5412
rect 4555 5468 4619 5472
rect 4555 5412 4559 5468
rect 4559 5412 4615 5468
rect 4615 5412 4619 5468
rect 4555 5408 4619 5412
rect 4635 5468 4699 5472
rect 4635 5412 4639 5468
rect 4639 5412 4695 5468
rect 4695 5412 4699 5468
rect 4635 5408 4699 5412
rect 4715 5468 4779 5472
rect 4715 5412 4719 5468
rect 4719 5412 4775 5468
rect 4775 5412 4779 5468
rect 4715 5408 4779 5412
rect 10202 5468 10266 5472
rect 10202 5412 10206 5468
rect 10206 5412 10262 5468
rect 10262 5412 10266 5468
rect 10202 5408 10266 5412
rect 10282 5468 10346 5472
rect 10282 5412 10286 5468
rect 10286 5412 10342 5468
rect 10342 5412 10346 5468
rect 10282 5408 10346 5412
rect 10362 5468 10426 5472
rect 10362 5412 10366 5468
rect 10366 5412 10422 5468
rect 10422 5412 10426 5468
rect 10362 5408 10426 5412
rect 10442 5468 10506 5472
rect 10442 5412 10446 5468
rect 10446 5412 10502 5468
rect 10502 5412 10506 5468
rect 10442 5408 10506 5412
rect 15929 5468 15993 5472
rect 15929 5412 15933 5468
rect 15933 5412 15989 5468
rect 15989 5412 15993 5468
rect 15929 5408 15993 5412
rect 16009 5468 16073 5472
rect 16009 5412 16013 5468
rect 16013 5412 16069 5468
rect 16069 5412 16073 5468
rect 16009 5408 16073 5412
rect 16089 5468 16153 5472
rect 16089 5412 16093 5468
rect 16093 5412 16149 5468
rect 16149 5412 16153 5468
rect 16089 5408 16153 5412
rect 16169 5468 16233 5472
rect 16169 5412 16173 5468
rect 16173 5412 16229 5468
rect 16229 5412 16233 5468
rect 16169 5408 16233 5412
rect 21656 5468 21720 5472
rect 21656 5412 21660 5468
rect 21660 5412 21716 5468
rect 21716 5412 21720 5468
rect 21656 5408 21720 5412
rect 21736 5468 21800 5472
rect 21736 5412 21740 5468
rect 21740 5412 21796 5468
rect 21796 5412 21800 5468
rect 21736 5408 21800 5412
rect 21816 5468 21880 5472
rect 21816 5412 21820 5468
rect 21820 5412 21876 5468
rect 21876 5412 21880 5468
rect 21816 5408 21880 5412
rect 21896 5468 21960 5472
rect 21896 5412 21900 5468
rect 21900 5412 21956 5468
rect 21956 5412 21960 5468
rect 21896 5408 21960 5412
rect 3815 4924 3879 4928
rect 3815 4868 3819 4924
rect 3819 4868 3875 4924
rect 3875 4868 3879 4924
rect 3815 4864 3879 4868
rect 3895 4924 3959 4928
rect 3895 4868 3899 4924
rect 3899 4868 3955 4924
rect 3955 4868 3959 4924
rect 3895 4864 3959 4868
rect 3975 4924 4039 4928
rect 3975 4868 3979 4924
rect 3979 4868 4035 4924
rect 4035 4868 4039 4924
rect 3975 4864 4039 4868
rect 4055 4924 4119 4928
rect 4055 4868 4059 4924
rect 4059 4868 4115 4924
rect 4115 4868 4119 4924
rect 4055 4864 4119 4868
rect 9542 4924 9606 4928
rect 9542 4868 9546 4924
rect 9546 4868 9602 4924
rect 9602 4868 9606 4924
rect 9542 4864 9606 4868
rect 9622 4924 9686 4928
rect 9622 4868 9626 4924
rect 9626 4868 9682 4924
rect 9682 4868 9686 4924
rect 9622 4864 9686 4868
rect 9702 4924 9766 4928
rect 9702 4868 9706 4924
rect 9706 4868 9762 4924
rect 9762 4868 9766 4924
rect 9702 4864 9766 4868
rect 9782 4924 9846 4928
rect 9782 4868 9786 4924
rect 9786 4868 9842 4924
rect 9842 4868 9846 4924
rect 9782 4864 9846 4868
rect 15269 4924 15333 4928
rect 15269 4868 15273 4924
rect 15273 4868 15329 4924
rect 15329 4868 15333 4924
rect 15269 4864 15333 4868
rect 15349 4924 15413 4928
rect 15349 4868 15353 4924
rect 15353 4868 15409 4924
rect 15409 4868 15413 4924
rect 15349 4864 15413 4868
rect 15429 4924 15493 4928
rect 15429 4868 15433 4924
rect 15433 4868 15489 4924
rect 15489 4868 15493 4924
rect 15429 4864 15493 4868
rect 15509 4924 15573 4928
rect 15509 4868 15513 4924
rect 15513 4868 15569 4924
rect 15569 4868 15573 4924
rect 15509 4864 15573 4868
rect 20996 4924 21060 4928
rect 20996 4868 21000 4924
rect 21000 4868 21056 4924
rect 21056 4868 21060 4924
rect 20996 4864 21060 4868
rect 21076 4924 21140 4928
rect 21076 4868 21080 4924
rect 21080 4868 21136 4924
rect 21136 4868 21140 4924
rect 21076 4864 21140 4868
rect 21156 4924 21220 4928
rect 21156 4868 21160 4924
rect 21160 4868 21216 4924
rect 21216 4868 21220 4924
rect 21156 4864 21220 4868
rect 21236 4924 21300 4928
rect 21236 4868 21240 4924
rect 21240 4868 21296 4924
rect 21296 4868 21300 4924
rect 21236 4864 21300 4868
rect 4475 4380 4539 4384
rect 4475 4324 4479 4380
rect 4479 4324 4535 4380
rect 4535 4324 4539 4380
rect 4475 4320 4539 4324
rect 4555 4380 4619 4384
rect 4555 4324 4559 4380
rect 4559 4324 4615 4380
rect 4615 4324 4619 4380
rect 4555 4320 4619 4324
rect 4635 4380 4699 4384
rect 4635 4324 4639 4380
rect 4639 4324 4695 4380
rect 4695 4324 4699 4380
rect 4635 4320 4699 4324
rect 4715 4380 4779 4384
rect 4715 4324 4719 4380
rect 4719 4324 4775 4380
rect 4775 4324 4779 4380
rect 4715 4320 4779 4324
rect 10202 4380 10266 4384
rect 10202 4324 10206 4380
rect 10206 4324 10262 4380
rect 10262 4324 10266 4380
rect 10202 4320 10266 4324
rect 10282 4380 10346 4384
rect 10282 4324 10286 4380
rect 10286 4324 10342 4380
rect 10342 4324 10346 4380
rect 10282 4320 10346 4324
rect 10362 4380 10426 4384
rect 10362 4324 10366 4380
rect 10366 4324 10422 4380
rect 10422 4324 10426 4380
rect 10362 4320 10426 4324
rect 10442 4380 10506 4384
rect 10442 4324 10446 4380
rect 10446 4324 10502 4380
rect 10502 4324 10506 4380
rect 10442 4320 10506 4324
rect 15929 4380 15993 4384
rect 15929 4324 15933 4380
rect 15933 4324 15989 4380
rect 15989 4324 15993 4380
rect 15929 4320 15993 4324
rect 16009 4380 16073 4384
rect 16009 4324 16013 4380
rect 16013 4324 16069 4380
rect 16069 4324 16073 4380
rect 16009 4320 16073 4324
rect 16089 4380 16153 4384
rect 16089 4324 16093 4380
rect 16093 4324 16149 4380
rect 16149 4324 16153 4380
rect 16089 4320 16153 4324
rect 16169 4380 16233 4384
rect 16169 4324 16173 4380
rect 16173 4324 16229 4380
rect 16229 4324 16233 4380
rect 16169 4320 16233 4324
rect 21656 4380 21720 4384
rect 21656 4324 21660 4380
rect 21660 4324 21716 4380
rect 21716 4324 21720 4380
rect 21656 4320 21720 4324
rect 21736 4380 21800 4384
rect 21736 4324 21740 4380
rect 21740 4324 21796 4380
rect 21796 4324 21800 4380
rect 21736 4320 21800 4324
rect 21816 4380 21880 4384
rect 21816 4324 21820 4380
rect 21820 4324 21876 4380
rect 21876 4324 21880 4380
rect 21816 4320 21880 4324
rect 21896 4380 21960 4384
rect 21896 4324 21900 4380
rect 21900 4324 21956 4380
rect 21956 4324 21960 4380
rect 21896 4320 21960 4324
rect 3815 3836 3879 3840
rect 3815 3780 3819 3836
rect 3819 3780 3875 3836
rect 3875 3780 3879 3836
rect 3815 3776 3879 3780
rect 3895 3836 3959 3840
rect 3895 3780 3899 3836
rect 3899 3780 3955 3836
rect 3955 3780 3959 3836
rect 3895 3776 3959 3780
rect 3975 3836 4039 3840
rect 3975 3780 3979 3836
rect 3979 3780 4035 3836
rect 4035 3780 4039 3836
rect 3975 3776 4039 3780
rect 4055 3836 4119 3840
rect 4055 3780 4059 3836
rect 4059 3780 4115 3836
rect 4115 3780 4119 3836
rect 4055 3776 4119 3780
rect 9542 3836 9606 3840
rect 9542 3780 9546 3836
rect 9546 3780 9602 3836
rect 9602 3780 9606 3836
rect 9542 3776 9606 3780
rect 9622 3836 9686 3840
rect 9622 3780 9626 3836
rect 9626 3780 9682 3836
rect 9682 3780 9686 3836
rect 9622 3776 9686 3780
rect 9702 3836 9766 3840
rect 9702 3780 9706 3836
rect 9706 3780 9762 3836
rect 9762 3780 9766 3836
rect 9702 3776 9766 3780
rect 9782 3836 9846 3840
rect 9782 3780 9786 3836
rect 9786 3780 9842 3836
rect 9842 3780 9846 3836
rect 9782 3776 9846 3780
rect 15269 3836 15333 3840
rect 15269 3780 15273 3836
rect 15273 3780 15329 3836
rect 15329 3780 15333 3836
rect 15269 3776 15333 3780
rect 15349 3836 15413 3840
rect 15349 3780 15353 3836
rect 15353 3780 15409 3836
rect 15409 3780 15413 3836
rect 15349 3776 15413 3780
rect 15429 3836 15493 3840
rect 15429 3780 15433 3836
rect 15433 3780 15489 3836
rect 15489 3780 15493 3836
rect 15429 3776 15493 3780
rect 15509 3836 15573 3840
rect 15509 3780 15513 3836
rect 15513 3780 15569 3836
rect 15569 3780 15573 3836
rect 15509 3776 15573 3780
rect 20996 3836 21060 3840
rect 20996 3780 21000 3836
rect 21000 3780 21056 3836
rect 21056 3780 21060 3836
rect 20996 3776 21060 3780
rect 21076 3836 21140 3840
rect 21076 3780 21080 3836
rect 21080 3780 21136 3836
rect 21136 3780 21140 3836
rect 21076 3776 21140 3780
rect 21156 3836 21220 3840
rect 21156 3780 21160 3836
rect 21160 3780 21216 3836
rect 21216 3780 21220 3836
rect 21156 3776 21220 3780
rect 21236 3836 21300 3840
rect 21236 3780 21240 3836
rect 21240 3780 21296 3836
rect 21296 3780 21300 3836
rect 21236 3776 21300 3780
rect 4475 3292 4539 3296
rect 4475 3236 4479 3292
rect 4479 3236 4535 3292
rect 4535 3236 4539 3292
rect 4475 3232 4539 3236
rect 4555 3292 4619 3296
rect 4555 3236 4559 3292
rect 4559 3236 4615 3292
rect 4615 3236 4619 3292
rect 4555 3232 4619 3236
rect 4635 3292 4699 3296
rect 4635 3236 4639 3292
rect 4639 3236 4695 3292
rect 4695 3236 4699 3292
rect 4635 3232 4699 3236
rect 4715 3292 4779 3296
rect 4715 3236 4719 3292
rect 4719 3236 4775 3292
rect 4775 3236 4779 3292
rect 4715 3232 4779 3236
rect 10202 3292 10266 3296
rect 10202 3236 10206 3292
rect 10206 3236 10262 3292
rect 10262 3236 10266 3292
rect 10202 3232 10266 3236
rect 10282 3292 10346 3296
rect 10282 3236 10286 3292
rect 10286 3236 10342 3292
rect 10342 3236 10346 3292
rect 10282 3232 10346 3236
rect 10362 3292 10426 3296
rect 10362 3236 10366 3292
rect 10366 3236 10422 3292
rect 10422 3236 10426 3292
rect 10362 3232 10426 3236
rect 10442 3292 10506 3296
rect 10442 3236 10446 3292
rect 10446 3236 10502 3292
rect 10502 3236 10506 3292
rect 10442 3232 10506 3236
rect 15929 3292 15993 3296
rect 15929 3236 15933 3292
rect 15933 3236 15989 3292
rect 15989 3236 15993 3292
rect 15929 3232 15993 3236
rect 16009 3292 16073 3296
rect 16009 3236 16013 3292
rect 16013 3236 16069 3292
rect 16069 3236 16073 3292
rect 16009 3232 16073 3236
rect 16089 3292 16153 3296
rect 16089 3236 16093 3292
rect 16093 3236 16149 3292
rect 16149 3236 16153 3292
rect 16089 3232 16153 3236
rect 16169 3292 16233 3296
rect 16169 3236 16173 3292
rect 16173 3236 16229 3292
rect 16229 3236 16233 3292
rect 16169 3232 16233 3236
rect 21656 3292 21720 3296
rect 21656 3236 21660 3292
rect 21660 3236 21716 3292
rect 21716 3236 21720 3292
rect 21656 3232 21720 3236
rect 21736 3292 21800 3296
rect 21736 3236 21740 3292
rect 21740 3236 21796 3292
rect 21796 3236 21800 3292
rect 21736 3232 21800 3236
rect 21816 3292 21880 3296
rect 21816 3236 21820 3292
rect 21820 3236 21876 3292
rect 21876 3236 21880 3292
rect 21816 3232 21880 3236
rect 21896 3292 21960 3296
rect 21896 3236 21900 3292
rect 21900 3236 21956 3292
rect 21956 3236 21960 3292
rect 21896 3232 21960 3236
rect 3815 2748 3879 2752
rect 3815 2692 3819 2748
rect 3819 2692 3875 2748
rect 3875 2692 3879 2748
rect 3815 2688 3879 2692
rect 3895 2748 3959 2752
rect 3895 2692 3899 2748
rect 3899 2692 3955 2748
rect 3955 2692 3959 2748
rect 3895 2688 3959 2692
rect 3975 2748 4039 2752
rect 3975 2692 3979 2748
rect 3979 2692 4035 2748
rect 4035 2692 4039 2748
rect 3975 2688 4039 2692
rect 4055 2748 4119 2752
rect 4055 2692 4059 2748
rect 4059 2692 4115 2748
rect 4115 2692 4119 2748
rect 4055 2688 4119 2692
rect 9542 2748 9606 2752
rect 9542 2692 9546 2748
rect 9546 2692 9602 2748
rect 9602 2692 9606 2748
rect 9542 2688 9606 2692
rect 9622 2748 9686 2752
rect 9622 2692 9626 2748
rect 9626 2692 9682 2748
rect 9682 2692 9686 2748
rect 9622 2688 9686 2692
rect 9702 2748 9766 2752
rect 9702 2692 9706 2748
rect 9706 2692 9762 2748
rect 9762 2692 9766 2748
rect 9702 2688 9766 2692
rect 9782 2748 9846 2752
rect 9782 2692 9786 2748
rect 9786 2692 9842 2748
rect 9842 2692 9846 2748
rect 9782 2688 9846 2692
rect 15269 2748 15333 2752
rect 15269 2692 15273 2748
rect 15273 2692 15329 2748
rect 15329 2692 15333 2748
rect 15269 2688 15333 2692
rect 15349 2748 15413 2752
rect 15349 2692 15353 2748
rect 15353 2692 15409 2748
rect 15409 2692 15413 2748
rect 15349 2688 15413 2692
rect 15429 2748 15493 2752
rect 15429 2692 15433 2748
rect 15433 2692 15489 2748
rect 15489 2692 15493 2748
rect 15429 2688 15493 2692
rect 15509 2748 15573 2752
rect 15509 2692 15513 2748
rect 15513 2692 15569 2748
rect 15569 2692 15573 2748
rect 15509 2688 15573 2692
rect 20996 2748 21060 2752
rect 20996 2692 21000 2748
rect 21000 2692 21056 2748
rect 21056 2692 21060 2748
rect 20996 2688 21060 2692
rect 21076 2748 21140 2752
rect 21076 2692 21080 2748
rect 21080 2692 21136 2748
rect 21136 2692 21140 2748
rect 21076 2688 21140 2692
rect 21156 2748 21220 2752
rect 21156 2692 21160 2748
rect 21160 2692 21216 2748
rect 21216 2692 21220 2748
rect 21156 2688 21220 2692
rect 21236 2748 21300 2752
rect 21236 2692 21240 2748
rect 21240 2692 21296 2748
rect 21296 2692 21300 2748
rect 21236 2688 21300 2692
rect 4475 2204 4539 2208
rect 4475 2148 4479 2204
rect 4479 2148 4535 2204
rect 4535 2148 4539 2204
rect 4475 2144 4539 2148
rect 4555 2204 4619 2208
rect 4555 2148 4559 2204
rect 4559 2148 4615 2204
rect 4615 2148 4619 2204
rect 4555 2144 4619 2148
rect 4635 2204 4699 2208
rect 4635 2148 4639 2204
rect 4639 2148 4695 2204
rect 4695 2148 4699 2204
rect 4635 2144 4699 2148
rect 4715 2204 4779 2208
rect 4715 2148 4719 2204
rect 4719 2148 4775 2204
rect 4775 2148 4779 2204
rect 4715 2144 4779 2148
rect 10202 2204 10266 2208
rect 10202 2148 10206 2204
rect 10206 2148 10262 2204
rect 10262 2148 10266 2204
rect 10202 2144 10266 2148
rect 10282 2204 10346 2208
rect 10282 2148 10286 2204
rect 10286 2148 10342 2204
rect 10342 2148 10346 2204
rect 10282 2144 10346 2148
rect 10362 2204 10426 2208
rect 10362 2148 10366 2204
rect 10366 2148 10422 2204
rect 10422 2148 10426 2204
rect 10362 2144 10426 2148
rect 10442 2204 10506 2208
rect 10442 2148 10446 2204
rect 10446 2148 10502 2204
rect 10502 2148 10506 2204
rect 10442 2144 10506 2148
rect 15929 2204 15993 2208
rect 15929 2148 15933 2204
rect 15933 2148 15989 2204
rect 15989 2148 15993 2204
rect 15929 2144 15993 2148
rect 16009 2204 16073 2208
rect 16009 2148 16013 2204
rect 16013 2148 16069 2204
rect 16069 2148 16073 2204
rect 16009 2144 16073 2148
rect 16089 2204 16153 2208
rect 16089 2148 16093 2204
rect 16093 2148 16149 2204
rect 16149 2148 16153 2204
rect 16089 2144 16153 2148
rect 16169 2204 16233 2208
rect 16169 2148 16173 2204
rect 16173 2148 16229 2204
rect 16229 2148 16233 2204
rect 16169 2144 16233 2148
rect 21656 2204 21720 2208
rect 21656 2148 21660 2204
rect 21660 2148 21716 2204
rect 21716 2148 21720 2204
rect 21656 2144 21720 2148
rect 21736 2204 21800 2208
rect 21736 2148 21740 2204
rect 21740 2148 21796 2204
rect 21796 2148 21800 2204
rect 21736 2144 21800 2148
rect 21816 2204 21880 2208
rect 21816 2148 21820 2204
rect 21820 2148 21876 2204
rect 21876 2148 21880 2204
rect 21816 2144 21880 2148
rect 21896 2204 21960 2208
rect 21896 2148 21900 2204
rect 21900 2148 21956 2204
rect 21956 2148 21960 2204
rect 21896 2144 21960 2148
<< metal4 >>
rect 3807 24512 4127 25072
rect 3807 24448 3815 24512
rect 3879 24448 3895 24512
rect 3959 24448 3975 24512
rect 4039 24448 4055 24512
rect 4119 24448 4127 24512
rect 3807 23424 4127 24448
rect 3807 23360 3815 23424
rect 3879 23360 3895 23424
rect 3959 23360 3975 23424
rect 4039 23360 4055 23424
rect 4119 23360 4127 23424
rect 3807 22336 4127 23360
rect 3807 22272 3815 22336
rect 3879 22286 3895 22336
rect 3959 22286 3975 22336
rect 4039 22286 4055 22336
rect 4119 22272 4127 22336
rect 3807 22050 3849 22272
rect 4085 22050 4127 22272
rect 3807 21248 4127 22050
rect 3807 21184 3815 21248
rect 3879 21184 3895 21248
rect 3959 21184 3975 21248
rect 4039 21184 4055 21248
rect 4119 21184 4127 21248
rect 3807 20160 4127 21184
rect 3807 20096 3815 20160
rect 3879 20096 3895 20160
rect 3959 20096 3975 20160
rect 4039 20096 4055 20160
rect 4119 20096 4127 20160
rect 3807 19072 4127 20096
rect 3807 19008 3815 19072
rect 3879 19008 3895 19072
rect 3959 19008 3975 19072
rect 4039 19008 4055 19072
rect 4119 19008 4127 19072
rect 3807 17984 4127 19008
rect 3807 17920 3815 17984
rect 3879 17920 3895 17984
rect 3959 17920 3975 17984
rect 4039 17920 4055 17984
rect 4119 17920 4127 17984
rect 3807 16896 4127 17920
rect 3807 16832 3815 16896
rect 3879 16832 3895 16896
rect 3959 16832 3975 16896
rect 4039 16832 4055 16896
rect 4119 16832 4127 16896
rect 3807 16574 4127 16832
rect 3807 16338 3849 16574
rect 4085 16338 4127 16574
rect 3807 15808 4127 16338
rect 3807 15744 3815 15808
rect 3879 15744 3895 15808
rect 3959 15744 3975 15808
rect 4039 15744 4055 15808
rect 4119 15744 4127 15808
rect 3807 14720 4127 15744
rect 3807 14656 3815 14720
rect 3879 14656 3895 14720
rect 3959 14656 3975 14720
rect 4039 14656 4055 14720
rect 4119 14656 4127 14720
rect 3807 13632 4127 14656
rect 3807 13568 3815 13632
rect 3879 13568 3895 13632
rect 3959 13568 3975 13632
rect 4039 13568 4055 13632
rect 4119 13568 4127 13632
rect 3807 12544 4127 13568
rect 3807 12480 3815 12544
rect 3879 12480 3895 12544
rect 3959 12480 3975 12544
rect 4039 12480 4055 12544
rect 4119 12480 4127 12544
rect 3807 11456 4127 12480
rect 3807 11392 3815 11456
rect 3879 11392 3895 11456
rect 3959 11392 3975 11456
rect 4039 11392 4055 11456
rect 4119 11392 4127 11456
rect 3807 10862 4127 11392
rect 3807 10626 3849 10862
rect 4085 10626 4127 10862
rect 3807 10368 4127 10626
rect 3807 10304 3815 10368
rect 3879 10304 3895 10368
rect 3959 10304 3975 10368
rect 4039 10304 4055 10368
rect 4119 10304 4127 10368
rect 3807 9280 4127 10304
rect 3807 9216 3815 9280
rect 3879 9216 3895 9280
rect 3959 9216 3975 9280
rect 4039 9216 4055 9280
rect 4119 9216 4127 9280
rect 3807 8192 4127 9216
rect 3807 8128 3815 8192
rect 3879 8128 3895 8192
rect 3959 8128 3975 8192
rect 4039 8128 4055 8192
rect 4119 8128 4127 8192
rect 3807 7104 4127 8128
rect 3807 7040 3815 7104
rect 3879 7040 3895 7104
rect 3959 7040 3975 7104
rect 4039 7040 4055 7104
rect 4119 7040 4127 7104
rect 3807 6016 4127 7040
rect 3807 5952 3815 6016
rect 3879 5952 3895 6016
rect 3959 5952 3975 6016
rect 4039 5952 4055 6016
rect 4119 5952 4127 6016
rect 3807 5150 4127 5952
rect 3807 4928 3849 5150
rect 4085 4928 4127 5150
rect 3807 4864 3815 4928
rect 3879 4864 3895 4914
rect 3959 4864 3975 4914
rect 4039 4864 4055 4914
rect 4119 4864 4127 4928
rect 3807 3840 4127 4864
rect 3807 3776 3815 3840
rect 3879 3776 3895 3840
rect 3959 3776 3975 3840
rect 4039 3776 4055 3840
rect 4119 3776 4127 3840
rect 3807 2752 4127 3776
rect 3807 2688 3815 2752
rect 3879 2688 3895 2752
rect 3959 2688 3975 2752
rect 4039 2688 4055 2752
rect 4119 2688 4127 2752
rect 3807 2128 4127 2688
rect 4467 25056 4787 25072
rect 4467 24992 4475 25056
rect 4539 24992 4555 25056
rect 4619 24992 4635 25056
rect 4699 24992 4715 25056
rect 4779 24992 4787 25056
rect 4467 23968 4787 24992
rect 4467 23904 4475 23968
rect 4539 23904 4555 23968
rect 4619 23904 4635 23968
rect 4699 23904 4715 23968
rect 4779 23904 4787 23968
rect 4467 22946 4787 23904
rect 4467 22880 4509 22946
rect 4745 22880 4787 22946
rect 4467 22816 4475 22880
rect 4779 22816 4787 22880
rect 4467 22710 4509 22816
rect 4745 22710 4787 22816
rect 4467 21792 4787 22710
rect 4467 21728 4475 21792
rect 4539 21728 4555 21792
rect 4619 21728 4635 21792
rect 4699 21728 4715 21792
rect 4779 21728 4787 21792
rect 4467 20704 4787 21728
rect 4467 20640 4475 20704
rect 4539 20640 4555 20704
rect 4619 20640 4635 20704
rect 4699 20640 4715 20704
rect 4779 20640 4787 20704
rect 4467 19616 4787 20640
rect 4467 19552 4475 19616
rect 4539 19552 4555 19616
rect 4619 19552 4635 19616
rect 4699 19552 4715 19616
rect 4779 19552 4787 19616
rect 4467 18528 4787 19552
rect 4467 18464 4475 18528
rect 4539 18464 4555 18528
rect 4619 18464 4635 18528
rect 4699 18464 4715 18528
rect 4779 18464 4787 18528
rect 4467 17440 4787 18464
rect 4467 17376 4475 17440
rect 4539 17376 4555 17440
rect 4619 17376 4635 17440
rect 4699 17376 4715 17440
rect 4779 17376 4787 17440
rect 4467 17234 4787 17376
rect 4467 16998 4509 17234
rect 4745 16998 4787 17234
rect 4467 16352 4787 16998
rect 4467 16288 4475 16352
rect 4539 16288 4555 16352
rect 4619 16288 4635 16352
rect 4699 16288 4715 16352
rect 4779 16288 4787 16352
rect 4467 15264 4787 16288
rect 4467 15200 4475 15264
rect 4539 15200 4555 15264
rect 4619 15200 4635 15264
rect 4699 15200 4715 15264
rect 4779 15200 4787 15264
rect 4467 14176 4787 15200
rect 4467 14112 4475 14176
rect 4539 14112 4555 14176
rect 4619 14112 4635 14176
rect 4699 14112 4715 14176
rect 4779 14112 4787 14176
rect 4467 13088 4787 14112
rect 4467 13024 4475 13088
rect 4539 13024 4555 13088
rect 4619 13024 4635 13088
rect 4699 13024 4715 13088
rect 4779 13024 4787 13088
rect 4467 12000 4787 13024
rect 4467 11936 4475 12000
rect 4539 11936 4555 12000
rect 4619 11936 4635 12000
rect 4699 11936 4715 12000
rect 4779 11936 4787 12000
rect 4467 11522 4787 11936
rect 4467 11286 4509 11522
rect 4745 11286 4787 11522
rect 4467 10912 4787 11286
rect 4467 10848 4475 10912
rect 4539 10848 4555 10912
rect 4619 10848 4635 10912
rect 4699 10848 4715 10912
rect 4779 10848 4787 10912
rect 4467 9824 4787 10848
rect 4467 9760 4475 9824
rect 4539 9760 4555 9824
rect 4619 9760 4635 9824
rect 4699 9760 4715 9824
rect 4779 9760 4787 9824
rect 4467 8736 4787 9760
rect 4467 8672 4475 8736
rect 4539 8672 4555 8736
rect 4619 8672 4635 8736
rect 4699 8672 4715 8736
rect 4779 8672 4787 8736
rect 4467 7648 4787 8672
rect 4467 7584 4475 7648
rect 4539 7584 4555 7648
rect 4619 7584 4635 7648
rect 4699 7584 4715 7648
rect 4779 7584 4787 7648
rect 4467 6560 4787 7584
rect 4467 6496 4475 6560
rect 4539 6496 4555 6560
rect 4619 6496 4635 6560
rect 4699 6496 4715 6560
rect 4779 6496 4787 6560
rect 4467 5810 4787 6496
rect 4467 5574 4509 5810
rect 4745 5574 4787 5810
rect 4467 5472 4787 5574
rect 4467 5408 4475 5472
rect 4539 5408 4555 5472
rect 4619 5408 4635 5472
rect 4699 5408 4715 5472
rect 4779 5408 4787 5472
rect 4467 4384 4787 5408
rect 4467 4320 4475 4384
rect 4539 4320 4555 4384
rect 4619 4320 4635 4384
rect 4699 4320 4715 4384
rect 4779 4320 4787 4384
rect 4467 3296 4787 4320
rect 4467 3232 4475 3296
rect 4539 3232 4555 3296
rect 4619 3232 4635 3296
rect 4699 3232 4715 3296
rect 4779 3232 4787 3296
rect 4467 2208 4787 3232
rect 4467 2144 4475 2208
rect 4539 2144 4555 2208
rect 4619 2144 4635 2208
rect 4699 2144 4715 2208
rect 4779 2144 4787 2208
rect 4467 2128 4787 2144
rect 9534 24512 9854 25072
rect 9534 24448 9542 24512
rect 9606 24448 9622 24512
rect 9686 24448 9702 24512
rect 9766 24448 9782 24512
rect 9846 24448 9854 24512
rect 9534 23424 9854 24448
rect 9534 23360 9542 23424
rect 9606 23360 9622 23424
rect 9686 23360 9702 23424
rect 9766 23360 9782 23424
rect 9846 23360 9854 23424
rect 9534 22336 9854 23360
rect 9534 22272 9542 22336
rect 9606 22286 9622 22336
rect 9686 22286 9702 22336
rect 9766 22286 9782 22336
rect 9846 22272 9854 22336
rect 9534 22050 9576 22272
rect 9812 22050 9854 22272
rect 9534 21248 9854 22050
rect 9534 21184 9542 21248
rect 9606 21184 9622 21248
rect 9686 21184 9702 21248
rect 9766 21184 9782 21248
rect 9846 21184 9854 21248
rect 9534 20160 9854 21184
rect 9534 20096 9542 20160
rect 9606 20096 9622 20160
rect 9686 20096 9702 20160
rect 9766 20096 9782 20160
rect 9846 20096 9854 20160
rect 9534 19072 9854 20096
rect 9534 19008 9542 19072
rect 9606 19008 9622 19072
rect 9686 19008 9702 19072
rect 9766 19008 9782 19072
rect 9846 19008 9854 19072
rect 9534 17984 9854 19008
rect 9534 17920 9542 17984
rect 9606 17920 9622 17984
rect 9686 17920 9702 17984
rect 9766 17920 9782 17984
rect 9846 17920 9854 17984
rect 9534 16896 9854 17920
rect 9534 16832 9542 16896
rect 9606 16832 9622 16896
rect 9686 16832 9702 16896
rect 9766 16832 9782 16896
rect 9846 16832 9854 16896
rect 9534 16574 9854 16832
rect 9534 16338 9576 16574
rect 9812 16338 9854 16574
rect 9534 15808 9854 16338
rect 9534 15744 9542 15808
rect 9606 15744 9622 15808
rect 9686 15744 9702 15808
rect 9766 15744 9782 15808
rect 9846 15744 9854 15808
rect 9534 14720 9854 15744
rect 9534 14656 9542 14720
rect 9606 14656 9622 14720
rect 9686 14656 9702 14720
rect 9766 14656 9782 14720
rect 9846 14656 9854 14720
rect 9534 13632 9854 14656
rect 9534 13568 9542 13632
rect 9606 13568 9622 13632
rect 9686 13568 9702 13632
rect 9766 13568 9782 13632
rect 9846 13568 9854 13632
rect 9534 12544 9854 13568
rect 9534 12480 9542 12544
rect 9606 12480 9622 12544
rect 9686 12480 9702 12544
rect 9766 12480 9782 12544
rect 9846 12480 9854 12544
rect 9534 11456 9854 12480
rect 9534 11392 9542 11456
rect 9606 11392 9622 11456
rect 9686 11392 9702 11456
rect 9766 11392 9782 11456
rect 9846 11392 9854 11456
rect 9534 10862 9854 11392
rect 9534 10626 9576 10862
rect 9812 10626 9854 10862
rect 9534 10368 9854 10626
rect 9534 10304 9542 10368
rect 9606 10304 9622 10368
rect 9686 10304 9702 10368
rect 9766 10304 9782 10368
rect 9846 10304 9854 10368
rect 9534 9280 9854 10304
rect 9534 9216 9542 9280
rect 9606 9216 9622 9280
rect 9686 9216 9702 9280
rect 9766 9216 9782 9280
rect 9846 9216 9854 9280
rect 9534 8192 9854 9216
rect 9534 8128 9542 8192
rect 9606 8128 9622 8192
rect 9686 8128 9702 8192
rect 9766 8128 9782 8192
rect 9846 8128 9854 8192
rect 9534 7104 9854 8128
rect 9534 7040 9542 7104
rect 9606 7040 9622 7104
rect 9686 7040 9702 7104
rect 9766 7040 9782 7104
rect 9846 7040 9854 7104
rect 9534 6016 9854 7040
rect 9534 5952 9542 6016
rect 9606 5952 9622 6016
rect 9686 5952 9702 6016
rect 9766 5952 9782 6016
rect 9846 5952 9854 6016
rect 9534 5150 9854 5952
rect 9534 4928 9576 5150
rect 9812 4928 9854 5150
rect 9534 4864 9542 4928
rect 9606 4864 9622 4914
rect 9686 4864 9702 4914
rect 9766 4864 9782 4914
rect 9846 4864 9854 4928
rect 9534 3840 9854 4864
rect 9534 3776 9542 3840
rect 9606 3776 9622 3840
rect 9686 3776 9702 3840
rect 9766 3776 9782 3840
rect 9846 3776 9854 3840
rect 9534 2752 9854 3776
rect 9534 2688 9542 2752
rect 9606 2688 9622 2752
rect 9686 2688 9702 2752
rect 9766 2688 9782 2752
rect 9846 2688 9854 2752
rect 9534 2128 9854 2688
rect 10194 25056 10514 25072
rect 10194 24992 10202 25056
rect 10266 24992 10282 25056
rect 10346 24992 10362 25056
rect 10426 24992 10442 25056
rect 10506 24992 10514 25056
rect 10194 23968 10514 24992
rect 10194 23904 10202 23968
rect 10266 23904 10282 23968
rect 10346 23904 10362 23968
rect 10426 23904 10442 23968
rect 10506 23904 10514 23968
rect 10194 22946 10514 23904
rect 10194 22880 10236 22946
rect 10472 22880 10514 22946
rect 10194 22816 10202 22880
rect 10506 22816 10514 22880
rect 10194 22710 10236 22816
rect 10472 22710 10514 22816
rect 10194 21792 10514 22710
rect 10194 21728 10202 21792
rect 10266 21728 10282 21792
rect 10346 21728 10362 21792
rect 10426 21728 10442 21792
rect 10506 21728 10514 21792
rect 10194 20704 10514 21728
rect 10194 20640 10202 20704
rect 10266 20640 10282 20704
rect 10346 20640 10362 20704
rect 10426 20640 10442 20704
rect 10506 20640 10514 20704
rect 10194 19616 10514 20640
rect 10194 19552 10202 19616
rect 10266 19552 10282 19616
rect 10346 19552 10362 19616
rect 10426 19552 10442 19616
rect 10506 19552 10514 19616
rect 10194 18528 10514 19552
rect 10194 18464 10202 18528
rect 10266 18464 10282 18528
rect 10346 18464 10362 18528
rect 10426 18464 10442 18528
rect 10506 18464 10514 18528
rect 10194 17440 10514 18464
rect 10194 17376 10202 17440
rect 10266 17376 10282 17440
rect 10346 17376 10362 17440
rect 10426 17376 10442 17440
rect 10506 17376 10514 17440
rect 10194 17234 10514 17376
rect 10194 16998 10236 17234
rect 10472 16998 10514 17234
rect 10194 16352 10514 16998
rect 10194 16288 10202 16352
rect 10266 16288 10282 16352
rect 10346 16288 10362 16352
rect 10426 16288 10442 16352
rect 10506 16288 10514 16352
rect 10194 15264 10514 16288
rect 10194 15200 10202 15264
rect 10266 15200 10282 15264
rect 10346 15200 10362 15264
rect 10426 15200 10442 15264
rect 10506 15200 10514 15264
rect 10194 14176 10514 15200
rect 10194 14112 10202 14176
rect 10266 14112 10282 14176
rect 10346 14112 10362 14176
rect 10426 14112 10442 14176
rect 10506 14112 10514 14176
rect 10194 13088 10514 14112
rect 10194 13024 10202 13088
rect 10266 13024 10282 13088
rect 10346 13024 10362 13088
rect 10426 13024 10442 13088
rect 10506 13024 10514 13088
rect 10194 12000 10514 13024
rect 10194 11936 10202 12000
rect 10266 11936 10282 12000
rect 10346 11936 10362 12000
rect 10426 11936 10442 12000
rect 10506 11936 10514 12000
rect 10194 11522 10514 11936
rect 10194 11286 10236 11522
rect 10472 11286 10514 11522
rect 10194 10912 10514 11286
rect 10194 10848 10202 10912
rect 10266 10848 10282 10912
rect 10346 10848 10362 10912
rect 10426 10848 10442 10912
rect 10506 10848 10514 10912
rect 10194 9824 10514 10848
rect 10194 9760 10202 9824
rect 10266 9760 10282 9824
rect 10346 9760 10362 9824
rect 10426 9760 10442 9824
rect 10506 9760 10514 9824
rect 10194 8736 10514 9760
rect 10194 8672 10202 8736
rect 10266 8672 10282 8736
rect 10346 8672 10362 8736
rect 10426 8672 10442 8736
rect 10506 8672 10514 8736
rect 10194 7648 10514 8672
rect 10194 7584 10202 7648
rect 10266 7584 10282 7648
rect 10346 7584 10362 7648
rect 10426 7584 10442 7648
rect 10506 7584 10514 7648
rect 10194 6560 10514 7584
rect 10194 6496 10202 6560
rect 10266 6496 10282 6560
rect 10346 6496 10362 6560
rect 10426 6496 10442 6560
rect 10506 6496 10514 6560
rect 10194 5810 10514 6496
rect 10194 5574 10236 5810
rect 10472 5574 10514 5810
rect 10194 5472 10514 5574
rect 10194 5408 10202 5472
rect 10266 5408 10282 5472
rect 10346 5408 10362 5472
rect 10426 5408 10442 5472
rect 10506 5408 10514 5472
rect 10194 4384 10514 5408
rect 10194 4320 10202 4384
rect 10266 4320 10282 4384
rect 10346 4320 10362 4384
rect 10426 4320 10442 4384
rect 10506 4320 10514 4384
rect 10194 3296 10514 4320
rect 10194 3232 10202 3296
rect 10266 3232 10282 3296
rect 10346 3232 10362 3296
rect 10426 3232 10442 3296
rect 10506 3232 10514 3296
rect 10194 2208 10514 3232
rect 10194 2144 10202 2208
rect 10266 2144 10282 2208
rect 10346 2144 10362 2208
rect 10426 2144 10442 2208
rect 10506 2144 10514 2208
rect 10194 2128 10514 2144
rect 15261 24512 15581 25072
rect 15261 24448 15269 24512
rect 15333 24448 15349 24512
rect 15413 24448 15429 24512
rect 15493 24448 15509 24512
rect 15573 24448 15581 24512
rect 15261 23424 15581 24448
rect 15261 23360 15269 23424
rect 15333 23360 15349 23424
rect 15413 23360 15429 23424
rect 15493 23360 15509 23424
rect 15573 23360 15581 23424
rect 15261 22336 15581 23360
rect 15261 22272 15269 22336
rect 15333 22286 15349 22336
rect 15413 22286 15429 22336
rect 15493 22286 15509 22336
rect 15573 22272 15581 22336
rect 15261 22050 15303 22272
rect 15539 22050 15581 22272
rect 15261 21248 15581 22050
rect 15261 21184 15269 21248
rect 15333 21184 15349 21248
rect 15413 21184 15429 21248
rect 15493 21184 15509 21248
rect 15573 21184 15581 21248
rect 15261 20160 15581 21184
rect 15261 20096 15269 20160
rect 15333 20096 15349 20160
rect 15413 20096 15429 20160
rect 15493 20096 15509 20160
rect 15573 20096 15581 20160
rect 15261 19072 15581 20096
rect 15261 19008 15269 19072
rect 15333 19008 15349 19072
rect 15413 19008 15429 19072
rect 15493 19008 15509 19072
rect 15573 19008 15581 19072
rect 15261 17984 15581 19008
rect 15261 17920 15269 17984
rect 15333 17920 15349 17984
rect 15413 17920 15429 17984
rect 15493 17920 15509 17984
rect 15573 17920 15581 17984
rect 15261 16896 15581 17920
rect 15261 16832 15269 16896
rect 15333 16832 15349 16896
rect 15413 16832 15429 16896
rect 15493 16832 15509 16896
rect 15573 16832 15581 16896
rect 15261 16574 15581 16832
rect 15261 16338 15303 16574
rect 15539 16338 15581 16574
rect 15261 15808 15581 16338
rect 15261 15744 15269 15808
rect 15333 15744 15349 15808
rect 15413 15744 15429 15808
rect 15493 15744 15509 15808
rect 15573 15744 15581 15808
rect 15261 14720 15581 15744
rect 15261 14656 15269 14720
rect 15333 14656 15349 14720
rect 15413 14656 15429 14720
rect 15493 14656 15509 14720
rect 15573 14656 15581 14720
rect 15261 13632 15581 14656
rect 15261 13568 15269 13632
rect 15333 13568 15349 13632
rect 15413 13568 15429 13632
rect 15493 13568 15509 13632
rect 15573 13568 15581 13632
rect 15261 12544 15581 13568
rect 15261 12480 15269 12544
rect 15333 12480 15349 12544
rect 15413 12480 15429 12544
rect 15493 12480 15509 12544
rect 15573 12480 15581 12544
rect 15261 11456 15581 12480
rect 15261 11392 15269 11456
rect 15333 11392 15349 11456
rect 15413 11392 15429 11456
rect 15493 11392 15509 11456
rect 15573 11392 15581 11456
rect 15261 10862 15581 11392
rect 15261 10626 15303 10862
rect 15539 10626 15581 10862
rect 15261 10368 15581 10626
rect 15261 10304 15269 10368
rect 15333 10304 15349 10368
rect 15413 10304 15429 10368
rect 15493 10304 15509 10368
rect 15573 10304 15581 10368
rect 15261 9280 15581 10304
rect 15261 9216 15269 9280
rect 15333 9216 15349 9280
rect 15413 9216 15429 9280
rect 15493 9216 15509 9280
rect 15573 9216 15581 9280
rect 15261 8192 15581 9216
rect 15261 8128 15269 8192
rect 15333 8128 15349 8192
rect 15413 8128 15429 8192
rect 15493 8128 15509 8192
rect 15573 8128 15581 8192
rect 15261 7104 15581 8128
rect 15261 7040 15269 7104
rect 15333 7040 15349 7104
rect 15413 7040 15429 7104
rect 15493 7040 15509 7104
rect 15573 7040 15581 7104
rect 15261 6016 15581 7040
rect 15261 5952 15269 6016
rect 15333 5952 15349 6016
rect 15413 5952 15429 6016
rect 15493 5952 15509 6016
rect 15573 5952 15581 6016
rect 15261 5150 15581 5952
rect 15261 4928 15303 5150
rect 15539 4928 15581 5150
rect 15261 4864 15269 4928
rect 15333 4864 15349 4914
rect 15413 4864 15429 4914
rect 15493 4864 15509 4914
rect 15573 4864 15581 4928
rect 15261 3840 15581 4864
rect 15261 3776 15269 3840
rect 15333 3776 15349 3840
rect 15413 3776 15429 3840
rect 15493 3776 15509 3840
rect 15573 3776 15581 3840
rect 15261 2752 15581 3776
rect 15261 2688 15269 2752
rect 15333 2688 15349 2752
rect 15413 2688 15429 2752
rect 15493 2688 15509 2752
rect 15573 2688 15581 2752
rect 15261 2128 15581 2688
rect 15921 25056 16241 25072
rect 15921 24992 15929 25056
rect 15993 24992 16009 25056
rect 16073 24992 16089 25056
rect 16153 24992 16169 25056
rect 16233 24992 16241 25056
rect 15921 23968 16241 24992
rect 15921 23904 15929 23968
rect 15993 23904 16009 23968
rect 16073 23904 16089 23968
rect 16153 23904 16169 23968
rect 16233 23904 16241 23968
rect 15921 22946 16241 23904
rect 15921 22880 15963 22946
rect 16199 22880 16241 22946
rect 15921 22816 15929 22880
rect 16233 22816 16241 22880
rect 15921 22710 15963 22816
rect 16199 22710 16241 22816
rect 15921 21792 16241 22710
rect 15921 21728 15929 21792
rect 15993 21728 16009 21792
rect 16073 21728 16089 21792
rect 16153 21728 16169 21792
rect 16233 21728 16241 21792
rect 15921 20704 16241 21728
rect 15921 20640 15929 20704
rect 15993 20640 16009 20704
rect 16073 20640 16089 20704
rect 16153 20640 16169 20704
rect 16233 20640 16241 20704
rect 15921 19616 16241 20640
rect 15921 19552 15929 19616
rect 15993 19552 16009 19616
rect 16073 19552 16089 19616
rect 16153 19552 16169 19616
rect 16233 19552 16241 19616
rect 15921 18528 16241 19552
rect 15921 18464 15929 18528
rect 15993 18464 16009 18528
rect 16073 18464 16089 18528
rect 16153 18464 16169 18528
rect 16233 18464 16241 18528
rect 15921 17440 16241 18464
rect 15921 17376 15929 17440
rect 15993 17376 16009 17440
rect 16073 17376 16089 17440
rect 16153 17376 16169 17440
rect 16233 17376 16241 17440
rect 15921 17234 16241 17376
rect 15921 16998 15963 17234
rect 16199 16998 16241 17234
rect 15921 16352 16241 16998
rect 15921 16288 15929 16352
rect 15993 16288 16009 16352
rect 16073 16288 16089 16352
rect 16153 16288 16169 16352
rect 16233 16288 16241 16352
rect 15921 15264 16241 16288
rect 15921 15200 15929 15264
rect 15993 15200 16009 15264
rect 16073 15200 16089 15264
rect 16153 15200 16169 15264
rect 16233 15200 16241 15264
rect 15921 14176 16241 15200
rect 15921 14112 15929 14176
rect 15993 14112 16009 14176
rect 16073 14112 16089 14176
rect 16153 14112 16169 14176
rect 16233 14112 16241 14176
rect 15921 13088 16241 14112
rect 15921 13024 15929 13088
rect 15993 13024 16009 13088
rect 16073 13024 16089 13088
rect 16153 13024 16169 13088
rect 16233 13024 16241 13088
rect 15921 12000 16241 13024
rect 15921 11936 15929 12000
rect 15993 11936 16009 12000
rect 16073 11936 16089 12000
rect 16153 11936 16169 12000
rect 16233 11936 16241 12000
rect 15921 11522 16241 11936
rect 15921 11286 15963 11522
rect 16199 11286 16241 11522
rect 15921 10912 16241 11286
rect 15921 10848 15929 10912
rect 15993 10848 16009 10912
rect 16073 10848 16089 10912
rect 16153 10848 16169 10912
rect 16233 10848 16241 10912
rect 15921 9824 16241 10848
rect 15921 9760 15929 9824
rect 15993 9760 16009 9824
rect 16073 9760 16089 9824
rect 16153 9760 16169 9824
rect 16233 9760 16241 9824
rect 15921 8736 16241 9760
rect 15921 8672 15929 8736
rect 15993 8672 16009 8736
rect 16073 8672 16089 8736
rect 16153 8672 16169 8736
rect 16233 8672 16241 8736
rect 15921 7648 16241 8672
rect 15921 7584 15929 7648
rect 15993 7584 16009 7648
rect 16073 7584 16089 7648
rect 16153 7584 16169 7648
rect 16233 7584 16241 7648
rect 15921 6560 16241 7584
rect 15921 6496 15929 6560
rect 15993 6496 16009 6560
rect 16073 6496 16089 6560
rect 16153 6496 16169 6560
rect 16233 6496 16241 6560
rect 15921 5810 16241 6496
rect 15921 5574 15963 5810
rect 16199 5574 16241 5810
rect 15921 5472 16241 5574
rect 15921 5408 15929 5472
rect 15993 5408 16009 5472
rect 16073 5408 16089 5472
rect 16153 5408 16169 5472
rect 16233 5408 16241 5472
rect 15921 4384 16241 5408
rect 15921 4320 15929 4384
rect 15993 4320 16009 4384
rect 16073 4320 16089 4384
rect 16153 4320 16169 4384
rect 16233 4320 16241 4384
rect 15921 3296 16241 4320
rect 15921 3232 15929 3296
rect 15993 3232 16009 3296
rect 16073 3232 16089 3296
rect 16153 3232 16169 3296
rect 16233 3232 16241 3296
rect 15921 2208 16241 3232
rect 15921 2144 15929 2208
rect 15993 2144 16009 2208
rect 16073 2144 16089 2208
rect 16153 2144 16169 2208
rect 16233 2144 16241 2208
rect 15921 2128 16241 2144
rect 20988 24512 21308 25072
rect 20988 24448 20996 24512
rect 21060 24448 21076 24512
rect 21140 24448 21156 24512
rect 21220 24448 21236 24512
rect 21300 24448 21308 24512
rect 20988 23424 21308 24448
rect 20988 23360 20996 23424
rect 21060 23360 21076 23424
rect 21140 23360 21156 23424
rect 21220 23360 21236 23424
rect 21300 23360 21308 23424
rect 20988 22336 21308 23360
rect 20988 22272 20996 22336
rect 21060 22286 21076 22336
rect 21140 22286 21156 22336
rect 21220 22286 21236 22336
rect 21300 22272 21308 22336
rect 20988 22050 21030 22272
rect 21266 22050 21308 22272
rect 20988 21248 21308 22050
rect 20988 21184 20996 21248
rect 21060 21184 21076 21248
rect 21140 21184 21156 21248
rect 21220 21184 21236 21248
rect 21300 21184 21308 21248
rect 20988 20160 21308 21184
rect 20988 20096 20996 20160
rect 21060 20096 21076 20160
rect 21140 20096 21156 20160
rect 21220 20096 21236 20160
rect 21300 20096 21308 20160
rect 20988 19072 21308 20096
rect 20988 19008 20996 19072
rect 21060 19008 21076 19072
rect 21140 19008 21156 19072
rect 21220 19008 21236 19072
rect 21300 19008 21308 19072
rect 20988 17984 21308 19008
rect 20988 17920 20996 17984
rect 21060 17920 21076 17984
rect 21140 17920 21156 17984
rect 21220 17920 21236 17984
rect 21300 17920 21308 17984
rect 20988 16896 21308 17920
rect 20988 16832 20996 16896
rect 21060 16832 21076 16896
rect 21140 16832 21156 16896
rect 21220 16832 21236 16896
rect 21300 16832 21308 16896
rect 20988 16574 21308 16832
rect 20988 16338 21030 16574
rect 21266 16338 21308 16574
rect 20988 15808 21308 16338
rect 20988 15744 20996 15808
rect 21060 15744 21076 15808
rect 21140 15744 21156 15808
rect 21220 15744 21236 15808
rect 21300 15744 21308 15808
rect 20988 14720 21308 15744
rect 20988 14656 20996 14720
rect 21060 14656 21076 14720
rect 21140 14656 21156 14720
rect 21220 14656 21236 14720
rect 21300 14656 21308 14720
rect 20988 13632 21308 14656
rect 20988 13568 20996 13632
rect 21060 13568 21076 13632
rect 21140 13568 21156 13632
rect 21220 13568 21236 13632
rect 21300 13568 21308 13632
rect 20988 12544 21308 13568
rect 20988 12480 20996 12544
rect 21060 12480 21076 12544
rect 21140 12480 21156 12544
rect 21220 12480 21236 12544
rect 21300 12480 21308 12544
rect 20988 11456 21308 12480
rect 20988 11392 20996 11456
rect 21060 11392 21076 11456
rect 21140 11392 21156 11456
rect 21220 11392 21236 11456
rect 21300 11392 21308 11456
rect 20988 10862 21308 11392
rect 20988 10626 21030 10862
rect 21266 10626 21308 10862
rect 20988 10368 21308 10626
rect 20988 10304 20996 10368
rect 21060 10304 21076 10368
rect 21140 10304 21156 10368
rect 21220 10304 21236 10368
rect 21300 10304 21308 10368
rect 20988 9280 21308 10304
rect 20988 9216 20996 9280
rect 21060 9216 21076 9280
rect 21140 9216 21156 9280
rect 21220 9216 21236 9280
rect 21300 9216 21308 9280
rect 20988 8192 21308 9216
rect 20988 8128 20996 8192
rect 21060 8128 21076 8192
rect 21140 8128 21156 8192
rect 21220 8128 21236 8192
rect 21300 8128 21308 8192
rect 20988 7104 21308 8128
rect 20988 7040 20996 7104
rect 21060 7040 21076 7104
rect 21140 7040 21156 7104
rect 21220 7040 21236 7104
rect 21300 7040 21308 7104
rect 20988 6016 21308 7040
rect 20988 5952 20996 6016
rect 21060 5952 21076 6016
rect 21140 5952 21156 6016
rect 21220 5952 21236 6016
rect 21300 5952 21308 6016
rect 20988 5150 21308 5952
rect 20988 4928 21030 5150
rect 21266 4928 21308 5150
rect 20988 4864 20996 4928
rect 21060 4864 21076 4914
rect 21140 4864 21156 4914
rect 21220 4864 21236 4914
rect 21300 4864 21308 4928
rect 20988 3840 21308 4864
rect 20988 3776 20996 3840
rect 21060 3776 21076 3840
rect 21140 3776 21156 3840
rect 21220 3776 21236 3840
rect 21300 3776 21308 3840
rect 20988 2752 21308 3776
rect 20988 2688 20996 2752
rect 21060 2688 21076 2752
rect 21140 2688 21156 2752
rect 21220 2688 21236 2752
rect 21300 2688 21308 2752
rect 20988 2128 21308 2688
rect 21648 25056 21968 25072
rect 21648 24992 21656 25056
rect 21720 24992 21736 25056
rect 21800 24992 21816 25056
rect 21880 24992 21896 25056
rect 21960 24992 21968 25056
rect 21648 23968 21968 24992
rect 21648 23904 21656 23968
rect 21720 23904 21736 23968
rect 21800 23904 21816 23968
rect 21880 23904 21896 23968
rect 21960 23904 21968 23968
rect 21648 22946 21968 23904
rect 21648 22880 21690 22946
rect 21926 22880 21968 22946
rect 21648 22816 21656 22880
rect 21960 22816 21968 22880
rect 21648 22710 21690 22816
rect 21926 22710 21968 22816
rect 21648 21792 21968 22710
rect 21648 21728 21656 21792
rect 21720 21728 21736 21792
rect 21800 21728 21816 21792
rect 21880 21728 21896 21792
rect 21960 21728 21968 21792
rect 21648 20704 21968 21728
rect 21648 20640 21656 20704
rect 21720 20640 21736 20704
rect 21800 20640 21816 20704
rect 21880 20640 21896 20704
rect 21960 20640 21968 20704
rect 21648 19616 21968 20640
rect 21648 19552 21656 19616
rect 21720 19552 21736 19616
rect 21800 19552 21816 19616
rect 21880 19552 21896 19616
rect 21960 19552 21968 19616
rect 21648 18528 21968 19552
rect 21648 18464 21656 18528
rect 21720 18464 21736 18528
rect 21800 18464 21816 18528
rect 21880 18464 21896 18528
rect 21960 18464 21968 18528
rect 21648 17440 21968 18464
rect 21648 17376 21656 17440
rect 21720 17376 21736 17440
rect 21800 17376 21816 17440
rect 21880 17376 21896 17440
rect 21960 17376 21968 17440
rect 21648 17234 21968 17376
rect 21648 16998 21690 17234
rect 21926 16998 21968 17234
rect 21648 16352 21968 16998
rect 21648 16288 21656 16352
rect 21720 16288 21736 16352
rect 21800 16288 21816 16352
rect 21880 16288 21896 16352
rect 21960 16288 21968 16352
rect 21648 15264 21968 16288
rect 21648 15200 21656 15264
rect 21720 15200 21736 15264
rect 21800 15200 21816 15264
rect 21880 15200 21896 15264
rect 21960 15200 21968 15264
rect 21648 14176 21968 15200
rect 21648 14112 21656 14176
rect 21720 14112 21736 14176
rect 21800 14112 21816 14176
rect 21880 14112 21896 14176
rect 21960 14112 21968 14176
rect 21648 13088 21968 14112
rect 21648 13024 21656 13088
rect 21720 13024 21736 13088
rect 21800 13024 21816 13088
rect 21880 13024 21896 13088
rect 21960 13024 21968 13088
rect 21648 12000 21968 13024
rect 21648 11936 21656 12000
rect 21720 11936 21736 12000
rect 21800 11936 21816 12000
rect 21880 11936 21896 12000
rect 21960 11936 21968 12000
rect 21648 11522 21968 11936
rect 21648 11286 21690 11522
rect 21926 11286 21968 11522
rect 21648 10912 21968 11286
rect 21648 10848 21656 10912
rect 21720 10848 21736 10912
rect 21800 10848 21816 10912
rect 21880 10848 21896 10912
rect 21960 10848 21968 10912
rect 21648 9824 21968 10848
rect 21648 9760 21656 9824
rect 21720 9760 21736 9824
rect 21800 9760 21816 9824
rect 21880 9760 21896 9824
rect 21960 9760 21968 9824
rect 21648 8736 21968 9760
rect 21648 8672 21656 8736
rect 21720 8672 21736 8736
rect 21800 8672 21816 8736
rect 21880 8672 21896 8736
rect 21960 8672 21968 8736
rect 21648 7648 21968 8672
rect 21648 7584 21656 7648
rect 21720 7584 21736 7648
rect 21800 7584 21816 7648
rect 21880 7584 21896 7648
rect 21960 7584 21968 7648
rect 21648 6560 21968 7584
rect 21648 6496 21656 6560
rect 21720 6496 21736 6560
rect 21800 6496 21816 6560
rect 21880 6496 21896 6560
rect 21960 6496 21968 6560
rect 21648 5810 21968 6496
rect 21648 5574 21690 5810
rect 21926 5574 21968 5810
rect 21648 5472 21968 5574
rect 21648 5408 21656 5472
rect 21720 5408 21736 5472
rect 21800 5408 21816 5472
rect 21880 5408 21896 5472
rect 21960 5408 21968 5472
rect 21648 4384 21968 5408
rect 21648 4320 21656 4384
rect 21720 4320 21736 4384
rect 21800 4320 21816 4384
rect 21880 4320 21896 4384
rect 21960 4320 21968 4384
rect 21648 3296 21968 4320
rect 21648 3232 21656 3296
rect 21720 3232 21736 3296
rect 21800 3232 21816 3296
rect 21880 3232 21896 3296
rect 21960 3232 21968 3296
rect 21648 2208 21968 3232
rect 21648 2144 21656 2208
rect 21720 2144 21736 2208
rect 21800 2144 21816 2208
rect 21880 2144 21896 2208
rect 21960 2144 21968 2208
rect 21648 2128 21968 2144
<< via4 >>
rect 3849 22272 3879 22286
rect 3879 22272 3895 22286
rect 3895 22272 3959 22286
rect 3959 22272 3975 22286
rect 3975 22272 4039 22286
rect 4039 22272 4055 22286
rect 4055 22272 4085 22286
rect 3849 22050 4085 22272
rect 3849 16338 4085 16574
rect 3849 10626 4085 10862
rect 3849 4928 4085 5150
rect 3849 4914 3879 4928
rect 3879 4914 3895 4928
rect 3895 4914 3959 4928
rect 3959 4914 3975 4928
rect 3975 4914 4039 4928
rect 4039 4914 4055 4928
rect 4055 4914 4085 4928
rect 4509 22880 4745 22946
rect 4509 22816 4539 22880
rect 4539 22816 4555 22880
rect 4555 22816 4619 22880
rect 4619 22816 4635 22880
rect 4635 22816 4699 22880
rect 4699 22816 4715 22880
rect 4715 22816 4745 22880
rect 4509 22710 4745 22816
rect 4509 16998 4745 17234
rect 4509 11286 4745 11522
rect 4509 5574 4745 5810
rect 9576 22272 9606 22286
rect 9606 22272 9622 22286
rect 9622 22272 9686 22286
rect 9686 22272 9702 22286
rect 9702 22272 9766 22286
rect 9766 22272 9782 22286
rect 9782 22272 9812 22286
rect 9576 22050 9812 22272
rect 9576 16338 9812 16574
rect 9576 10626 9812 10862
rect 9576 4928 9812 5150
rect 9576 4914 9606 4928
rect 9606 4914 9622 4928
rect 9622 4914 9686 4928
rect 9686 4914 9702 4928
rect 9702 4914 9766 4928
rect 9766 4914 9782 4928
rect 9782 4914 9812 4928
rect 10236 22880 10472 22946
rect 10236 22816 10266 22880
rect 10266 22816 10282 22880
rect 10282 22816 10346 22880
rect 10346 22816 10362 22880
rect 10362 22816 10426 22880
rect 10426 22816 10442 22880
rect 10442 22816 10472 22880
rect 10236 22710 10472 22816
rect 10236 16998 10472 17234
rect 10236 11286 10472 11522
rect 10236 5574 10472 5810
rect 15303 22272 15333 22286
rect 15333 22272 15349 22286
rect 15349 22272 15413 22286
rect 15413 22272 15429 22286
rect 15429 22272 15493 22286
rect 15493 22272 15509 22286
rect 15509 22272 15539 22286
rect 15303 22050 15539 22272
rect 15303 16338 15539 16574
rect 15303 10626 15539 10862
rect 15303 4928 15539 5150
rect 15303 4914 15333 4928
rect 15333 4914 15349 4928
rect 15349 4914 15413 4928
rect 15413 4914 15429 4928
rect 15429 4914 15493 4928
rect 15493 4914 15509 4928
rect 15509 4914 15539 4928
rect 15963 22880 16199 22946
rect 15963 22816 15993 22880
rect 15993 22816 16009 22880
rect 16009 22816 16073 22880
rect 16073 22816 16089 22880
rect 16089 22816 16153 22880
rect 16153 22816 16169 22880
rect 16169 22816 16199 22880
rect 15963 22710 16199 22816
rect 15963 16998 16199 17234
rect 15963 11286 16199 11522
rect 15963 5574 16199 5810
rect 21030 22272 21060 22286
rect 21060 22272 21076 22286
rect 21076 22272 21140 22286
rect 21140 22272 21156 22286
rect 21156 22272 21220 22286
rect 21220 22272 21236 22286
rect 21236 22272 21266 22286
rect 21030 22050 21266 22272
rect 21030 16338 21266 16574
rect 21030 10626 21266 10862
rect 21030 4928 21266 5150
rect 21030 4914 21060 4928
rect 21060 4914 21076 4928
rect 21076 4914 21140 4928
rect 21140 4914 21156 4928
rect 21156 4914 21220 4928
rect 21220 4914 21236 4928
rect 21236 4914 21266 4928
rect 21690 22880 21926 22946
rect 21690 22816 21720 22880
rect 21720 22816 21736 22880
rect 21736 22816 21800 22880
rect 21800 22816 21816 22880
rect 21816 22816 21880 22880
rect 21880 22816 21896 22880
rect 21896 22816 21926 22880
rect 21690 22710 21926 22816
rect 21690 16998 21926 17234
rect 21690 11286 21926 11522
rect 21690 5574 21926 5810
<< metal5 >>
rect 1056 22946 24060 22988
rect 1056 22710 4509 22946
rect 4745 22710 10236 22946
rect 10472 22710 15963 22946
rect 16199 22710 21690 22946
rect 21926 22710 24060 22946
rect 1056 22668 24060 22710
rect 1056 22286 24060 22328
rect 1056 22050 3849 22286
rect 4085 22050 9576 22286
rect 9812 22050 15303 22286
rect 15539 22050 21030 22286
rect 21266 22050 24060 22286
rect 1056 22008 24060 22050
rect 1056 17234 24060 17276
rect 1056 16998 4509 17234
rect 4745 16998 10236 17234
rect 10472 16998 15963 17234
rect 16199 16998 21690 17234
rect 21926 16998 24060 17234
rect 1056 16956 24060 16998
rect 1056 16574 24060 16616
rect 1056 16338 3849 16574
rect 4085 16338 9576 16574
rect 9812 16338 15303 16574
rect 15539 16338 21030 16574
rect 21266 16338 24060 16574
rect 1056 16296 24060 16338
rect 1056 11522 24060 11564
rect 1056 11286 4509 11522
rect 4745 11286 10236 11522
rect 10472 11286 15963 11522
rect 16199 11286 21690 11522
rect 21926 11286 24060 11522
rect 1056 11244 24060 11286
rect 1056 10862 24060 10904
rect 1056 10626 3849 10862
rect 4085 10626 9576 10862
rect 9812 10626 15303 10862
rect 15539 10626 21030 10862
rect 21266 10626 24060 10862
rect 1056 10584 24060 10626
rect 1056 5810 24060 5852
rect 1056 5574 4509 5810
rect 4745 5574 10236 5810
rect 10472 5574 15963 5810
rect 16199 5574 21690 5810
rect 21926 5574 24060 5810
rect 1056 5532 24060 5574
rect 1056 5150 24060 5192
rect 1056 4914 3849 5150
rect 4085 4914 9576 5150
rect 9812 4914 15303 5150
rect 15539 4914 21030 5150
rect 21266 4914 24060 5150
rect 1056 4872 24060 4914
use sky130_fd_sc_hd__nor4_1  _1388_
timestamp 0
transform -1 0 18400 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1389_
timestamp 0
transform 1 0 17204 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1390_
timestamp 0
transform -1 0 9200 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1391_
timestamp 0
transform -1 0 9568 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _1392_
timestamp 0
transform 1 0 13156 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1393_
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1394_
timestamp 0
transform 1 0 15364 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1395_
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _1396_
timestamp 0
transform -1 0 6808 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _1397_
timestamp 0
transform 1 0 13616 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1398_
timestamp 0
transform -1 0 14352 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1399_
timestamp 0
transform 1 0 13892 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  _1400_
timestamp 0
transform -1 0 11500 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1401_
timestamp 0
transform -1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1402_
timestamp 0
transform -1 0 10028 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1403_
timestamp 0
transform -1 0 10396 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1404_
timestamp 0
transform -1 0 10304 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1405_
timestamp 0
transform -1 0 10580 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1406_
timestamp 0
transform 1 0 10212 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1407_
timestamp 0
transform -1 0 11316 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1408_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1409_
timestamp 0
transform 1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1410_
timestamp 0
transform 1 0 10304 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1411_
timestamp 0
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1412_
timestamp 0
transform 1 0 8004 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1413_
timestamp 0
transform 1 0 9108 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1414_
timestamp 0
transform 1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1415_
timestamp 0
transform -1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1416_
timestamp 0
transform 1 0 13524 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1417_
timestamp 0
transform 1 0 13064 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1418_
timestamp 0
transform -1 0 13524 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1419_
timestamp 0
transform -1 0 13800 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1420_
timestamp 0
transform 1 0 12696 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1421_
timestamp 0
transform -1 0 13984 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1422_
timestamp 0
transform -1 0 13892 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1423_
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1424_
timestamp 0
transform -1 0 13248 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1425__127
timestamp 0
transform -1 0 14168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1425_
timestamp 0
transform -1 0 13800 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1426_
timestamp 0
transform -1 0 13892 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1427_
timestamp 0
transform 1 0 13156 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1428_
timestamp 0
transform -1 0 5336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1429_
timestamp 0
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1430_
timestamp 0
transform 1 0 4324 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1431_
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1432_
timestamp 0
transform 1 0 3956 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1433_
timestamp 0
transform -1 0 3680 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1434_
timestamp 0
transform 1 0 3680 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1435_
timestamp 0
transform -1 0 5520 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1436_
timestamp 0
transform 1 0 4600 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1437_
timestamp 0
transform 1 0 4232 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1438_
timestamp 0
transform -1 0 3680 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1439__128
timestamp 0
transform -1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1439_
timestamp 0
transform 1 0 4784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1440_
timestamp 0
transform -1 0 5428 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1441_
timestamp 0
transform -1 0 5060 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1442_
timestamp 0
transform -1 0 4692 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1443_
timestamp 0
transform 1 0 3312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1444_
timestamp 0
transform 1 0 4324 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1445_
timestamp 0
transform -1 0 3864 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1446_
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1447_
timestamp 0
transform 1 0 3864 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1448_
timestamp 0
transform 1 0 3588 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1449_
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1450_
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1451_
timestamp 0
transform 1 0 3956 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1452_
timestamp 0
transform -1 0 4416 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1453__129
timestamp 0
transform -1 0 5336 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1453_
timestamp 0
transform 1 0 4232 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1454_
timestamp 0
transform -1 0 5060 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1455_
timestamp 0
transform -1 0 4876 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1456_
timestamp 0
transform -1 0 7452 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1457_
timestamp 0
transform -1 0 7544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1458_
timestamp 0
transform 1 0 6992 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1459_
timestamp 0
transform 1 0 6440 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1460_
timestamp 0
transform 1 0 7268 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1461_
timestamp 0
transform 1 0 6532 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1462_
timestamp 0
transform 1 0 5796 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1463_
timestamp 0
transform 1 0 6532 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1464_
timestamp 0
transform 1 0 6348 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1465_
timestamp 0
transform 1 0 6348 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1466_
timestamp 0
transform 1 0 6440 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1467__130
timestamp 0
transform -1 0 7268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 0
transform 1 0 6624 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1468_
timestamp 0
transform -1 0 7176 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1469_
timestamp 0
transform 1 0 6440 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1470_
timestamp 0
transform -1 0 10028 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1471_
timestamp 0
transform -1 0 9200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1472_
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1473_
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1474_
timestamp 0
transform -1 0 9936 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1475_
timestamp 0
transform 1 0 9844 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1476_
timestamp 0
transform 1 0 8372 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1477_
timestamp 0
transform 1 0 8924 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1478_
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1479_
timestamp 0
transform 1 0 8924 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1480_
timestamp 0
transform -1 0 8924 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1481__131
timestamp 0
transform -1 0 9844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1481_
timestamp 0
transform 1 0 8740 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1482_
timestamp 0
transform -1 0 9476 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1483_
timestamp 0
transform 1 0 9016 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1484_
timestamp 0
transform -1 0 13156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1485_
timestamp 0
transform -1 0 12788 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1486_
timestamp 0
transform -1 0 12144 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1487_
timestamp 0
transform -1 0 12604 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1488_
timestamp 0
transform -1 0 12328 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1489_
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1490_
timestamp 0
transform -1 0 11408 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1491_
timestamp 0
transform 1 0 12696 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1492_
timestamp 0
transform 1 0 10120 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 0
transform 1 0 12052 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1494_
timestamp 0
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1495__132
timestamp 0
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1495_
timestamp 0
transform 1 0 10120 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1496_
timestamp 0
transform 1 0 9292 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1497_
timestamp 0
transform 1 0 11408 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1498_
timestamp 0
transform -1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1499_
timestamp 0
transform -1 0 13156 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1500_
timestamp 0
transform -1 0 12880 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1501_
timestamp 0
transform -1 0 12420 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1502_
timestamp 0
transform 1 0 13064 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1503_
timestamp 0
transform 1 0 12696 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1504_
timestamp 0
transform 1 0 12052 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1505_
timestamp 0
transform 1 0 12972 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1506_
timestamp 0
transform -1 0 12972 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 0
transform 1 0 12420 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 0
transform 1 0 12328 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1509_
timestamp 0
transform 1 0 11500 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1509__133
timestamp 0
transform -1 0 12144 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1510_
timestamp 0
transform 1 0 10396 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1511_
timestamp 0
transform 1 0 11592 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1512_
timestamp 0
transform -1 0 16468 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1513_
timestamp 0
transform -1 0 16192 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1514_
timestamp 0
transform 1 0 15640 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1515_
timestamp 0
transform 1 0 15732 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1516_
timestamp 0
transform -1 0 15088 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1517_
timestamp 0
transform -1 0 15732 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1518_
timestamp 0
transform -1 0 15364 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1519_
timestamp 0
transform 1 0 14168 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1520_
timestamp 0
transform 1 0 14628 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 0
transform 1 0 15456 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 0
transform 1 0 15088 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1523__134
timestamp 0
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 0
transform -1 0 17756 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 0
transform -1 0 17020 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1526_
timestamp 0
transform 1 0 14720 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1527_
timestamp 0
transform -1 0 14904 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1528_
timestamp 0
transform 1 0 14260 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1529_
timestamp 0
transform -1 0 15180 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1530_
timestamp 0
transform 1 0 15272 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1531_
timestamp 0
transform 1 0 14536 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1532_
timestamp 0
transform -1 0 15640 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1533_
timestamp 0
transform 1 0 14720 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1534_
timestamp 0
transform 1 0 14352 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1535_
timestamp 0
transform 1 0 15088 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1536_
timestamp 0
transform 1 0 14260 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1537__135
timestamp 0
transform -1 0 15732 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1537_
timestamp 0
transform 1 0 14628 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1538_
timestamp 0
transform -1 0 14628 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1539_
timestamp 0
transform 1 0 14168 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1540_
timestamp 0
transform -1 0 18584 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1541_
timestamp 0
transform -1 0 18308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1542_
timestamp 0
transform 1 0 17020 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1543_
timestamp 0
transform -1 0 16836 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1544_
timestamp 0
transform 1 0 17848 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1545_
timestamp 0
transform 1 0 17296 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1546_
timestamp 0
transform -1 0 18308 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1547_
timestamp 0
transform 1 0 17388 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1548_
timestamp 0
transform 1 0 16744 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1549_
timestamp 0
transform 1 0 17388 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1550_
timestamp 0
transform 1 0 17204 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1551__105
timestamp 0
transform -1 0 17940 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 0
transform 1 0 16836 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1552_
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 0
transform 1 0 16836 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1554_
timestamp 0
transform -1 0 23184 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1555_
timestamp 0
transform -1 0 21160 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1556_
timestamp 0
transform 1 0 21068 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1557_
timestamp 0
transform -1 0 21436 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1558_
timestamp 0
transform 1 0 20516 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1559_
timestamp 0
transform -1 0 20976 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1560_
timestamp 0
transform -1 0 20516 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1561_
timestamp 0
transform 1 0 20056 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1562_
timestamp 0
transform 1 0 19412 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1563_
timestamp 0
transform 1 0 22080 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1564_
timestamp 0
transform 1 0 20056 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1565__106
timestamp 0
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1565_
timestamp 0
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1566_
timestamp 0
transform 1 0 18952 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 0
transform 1 0 20240 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1568_
timestamp 0
transform -1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1569_
timestamp 0
transform 1 0 10120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1570_
timestamp 0
transform -1 0 11132 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1571_
timestamp 0
transform -1 0 10304 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1572_
timestamp 0
transform -1 0 10764 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1573_
timestamp 0
transform 1 0 10948 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1574_
timestamp 0
transform 1 0 10304 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1575_
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1576_
timestamp 0
transform 1 0 10488 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1577_
timestamp 0
transform 1 0 11500 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1578_
timestamp 0
transform -1 0 10672 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1579__107
timestamp 0
transform -1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1579_
timestamp 0
transform 1 0 10488 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1580_
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1581_
timestamp 0
transform 1 0 10304 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1582_
timestamp 0
transform -1 0 23644 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1583_
timestamp 0
transform -1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1584_
timestamp 0
transform -1 0 22540 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1585_
timestamp 0
transform 1 0 22540 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1586_
timestamp 0
transform -1 0 21620 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1587_
timestamp 0
transform -1 0 22080 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1588_
timestamp 0
transform -1 0 22448 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1589_
timestamp 0
transform 1 0 20976 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1590_
timestamp 0
transform -1 0 20976 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1591_
timestamp 0
transform 1 0 22540 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1592_
timestamp 0
transform 1 0 22540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1593__108
timestamp 0
transform -1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1593_
timestamp 0
transform 1 0 19504 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1594_
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1595_
timestamp 0
transform 1 0 21344 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1596_
timestamp 0
transform -1 0 23644 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1597_
timestamp 0
transform -1 0 23644 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1598_
timestamp 0
transform -1 0 21252 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1599_
timestamp 0
transform -1 0 21896 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1600_
timestamp 0
transform -1 0 21712 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1601_
timestamp 0
transform -1 0 22356 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1602_
timestamp 0
transform -1 0 22448 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1603_
timestamp 0
transform -1 0 22264 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1604_
timestamp 0
transform -1 0 22448 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1605_
timestamp 0
transform 1 0 22540 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1606_
timestamp 0
transform 1 0 22540 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1607__109
timestamp 0
transform -1 0 20976 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1607_
timestamp 0
transform 1 0 20332 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1608_
timestamp 0
transform 1 0 19504 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1609_
timestamp 0
transform 1 0 20976 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1610_
timestamp 0
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1611_
timestamp 0
transform -1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1612_
timestamp 0
transform 1 0 17664 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1613_
timestamp 0
transform 1 0 18032 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1614_
timestamp 0
transform -1 0 17388 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1615_
timestamp 0
transform -1 0 17572 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1616_
timestamp 0
transform 1 0 17388 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1617_
timestamp 0
transform -1 0 18216 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1618_
timestamp 0
transform -1 0 19136 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1619_
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1620_
timestamp 0
transform -1 0 17664 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1621__110
timestamp 0
transform -1 0 19044 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 0
transform 1 0 18124 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1622_
timestamp 0
transform -1 0 18492 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1623_
timestamp 0
transform -1 0 18492 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1624_
timestamp 0
transform -1 0 14720 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1625_
timestamp 0
transform -1 0 14352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1626_
timestamp 0
transform 1 0 13800 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1627_
timestamp 0
transform 1 0 13524 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1628_
timestamp 0
transform 1 0 15272 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1629_
timestamp 0
transform 1 0 14352 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1630_
timestamp 0
transform 1 0 14260 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1631_
timestamp 0
transform -1 0 15732 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1632_
timestamp 0
transform -1 0 15732 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1633_
timestamp 0
transform -1 0 14444 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1634_
timestamp 0
transform -1 0 13892 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1635__111
timestamp 0
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1635_
timestamp 0
transform 1 0 14904 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1636_
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1637_
timestamp 0
transform -1 0 14904 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1638_
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1639_
timestamp 0
transform -1 0 15272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1640_
timestamp 0
transform 1 0 15732 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1641_
timestamp 0
transform 1 0 15272 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1642_
timestamp 0
transform 1 0 16468 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1643_
timestamp 0
transform 1 0 15640 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1644_
timestamp 0
transform 1 0 15364 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1645_
timestamp 0
transform 1 0 16008 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1646_
timestamp 0
transform 1 0 15640 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1648_
timestamp 0
transform -1 0 14996 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1649__112
timestamp 0
transform -1 0 16468 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1649_
timestamp 0
transform 1 0 15732 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 0
transform -1 0 16100 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1651_
timestamp 0
transform 1 0 15364 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1652_
timestamp 0
transform -1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1653_
timestamp 0
transform -1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1654_
timestamp 0
transform -1 0 19688 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1655_
timestamp 0
transform -1 0 20056 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1656_
timestamp 0
transform -1 0 20240 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1657_
timestamp 0
transform 1 0 19872 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1658_
timestamp 0
transform -1 0 19872 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1659_
timestamp 0
transform 1 0 18768 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1660_
timestamp 0
transform -1 0 18768 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1661_
timestamp 0
transform 1 0 20424 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1662_
timestamp 0
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1663__113
timestamp 0
transform -1 0 18952 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1663_
timestamp 0
transform 1 0 18032 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1664_
timestamp 0
transform 1 0 17848 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 0
transform 1 0 18768 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1666_
timestamp 0
transform -1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1667_
timestamp 0
transform -1 0 23736 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1668_
timestamp 0
transform -1 0 22540 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1669_
timestamp 0
transform 1 0 21620 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1670_
timestamp 0
transform -1 0 21712 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1671_
timestamp 0
transform -1 0 22172 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1672_
timestamp 0
transform -1 0 21712 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1673_
timestamp 0
transform 1 0 20884 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1674_
timestamp 0
transform -1 0 20976 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 0
transform 1 0 22540 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1676_
timestamp 0
transform 1 0 22632 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1677__114
timestamp 0
transform 1 0 19780 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 0
transform 1 0 20056 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1680_
timestamp 0
transform -1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1681_
timestamp 0
transform -1 0 23092 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1682_
timestamp 0
transform -1 0 22724 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1683_
timestamp 0
transform -1 0 22264 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1684_
timestamp 0
transform -1 0 21804 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1685_
timestamp 0
transform -1 0 22264 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1686_
timestamp 0
transform -1 0 22448 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1687_
timestamp 0
transform 1 0 22080 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1688_
timestamp 0
transform -1 0 21712 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 0
transform 1 0 22540 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 0
transform 1 0 22540 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1691__115
timestamp 0
transform -1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1691_
timestamp 0
transform 1 0 20424 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1692_
timestamp 0
transform 1 0 19504 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1693_
timestamp 0
transform 1 0 21252 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1694_
timestamp 0
transform 1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1695_
timestamp 0
transform -1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1696_
timestamp 0
transform -1 0 19136 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1697_
timestamp 0
transform -1 0 20148 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1698_
timestamp 0
transform -1 0 18768 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1699_
timestamp 0
transform -1 0 19688 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1700_
timestamp 0
transform -1 0 20240 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1701_
timestamp 0
transform -1 0 19136 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1702_
timestamp 0
transform 1 0 18492 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 0
transform 1 0 20700 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1704_
timestamp 0
transform 1 0 19872 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1705__116
timestamp 0
transform -1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 0
transform 1 0 18676 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1706_
timestamp 0
transform 1 0 17848 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1707_
timestamp 0
transform 1 0 18768 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1708_
timestamp 0
transform -1 0 19044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1709_
timestamp 0
transform -1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1710_
timestamp 0
transform -1 0 17296 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1711_
timestamp 0
transform -1 0 18216 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1712_
timestamp 0
transform 1 0 17848 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1713_
timestamp 0
transform 1 0 17296 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1714_
timestamp 0
transform -1 0 18676 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1715_
timestamp 0
transform 1 0 17388 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1716_
timestamp 0
transform -1 0 17848 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 0
transform 1 0 18308 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1718_
timestamp 0
transform 1 0 17664 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1719__117
timestamp 0
transform -1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1719_
timestamp 0
transform 1 0 17112 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1720_
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1721_
timestamp 0
transform 1 0 17204 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1722_
timestamp 0
transform -1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1723_
timestamp 0
transform -1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1724_
timestamp 0
transform 1 0 7912 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1725_
timestamp 0
transform 1 0 7544 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1726_
timestamp 0
transform 1 0 7452 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1727_
timestamp 0
transform 1 0 6624 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1728_
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1729_
timestamp 0
transform -1 0 9016 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1730_
timestamp 0
transform 1 0 7912 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1731_
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1732_
timestamp 0
transform 1 0 6624 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1733__118
timestamp 0
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 0
transform 1 0 8648 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1734_
timestamp 0
transform -1 0 8648 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1735_
timestamp 0
transform -1 0 8556 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1736_
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1737_
timestamp 0
transform -1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1738_
timestamp 0
transform 1 0 15640 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1739_
timestamp 0
transform 1 0 14812 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1740_
timestamp 0
transform -1 0 14812 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1741_
timestamp 0
transform 1 0 14352 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1742_
timestamp 0
transform 1 0 14168 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1743_
timestamp 0
transform -1 0 15364 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1744_
timestamp 0
transform 1 0 15180 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1745_
timestamp 0
transform 1 0 15456 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 0
transform 1 0 14628 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1747__119
timestamp 0
transform -1 0 16468 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1747_
timestamp 0
transform 1 0 15364 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 0
transform 1 0 14996 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1749_
timestamp 0
transform -1 0 15640 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1750_
timestamp 0
transform -1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1751_
timestamp 0
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1752_
timestamp 0
transform -1 0 4140 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1753_
timestamp 0
transform 1 0 4600 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1754_
timestamp 0
transform 1 0 4600 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1755_
timestamp 0
transform 1 0 4140 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1756_
timestamp 0
transform 1 0 4600 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1757_
timestamp 0
transform -1 0 5704 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1758_
timestamp 0
transform -1 0 6164 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 0
transform 1 0 4784 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1760_
timestamp 0
transform 1 0 4600 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1761__120
timestamp 0
transform -1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1762_
timestamp 0
transform -1 0 5612 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 0
transform -1 0 5520 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1764_
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1765_
timestamp 0
transform 1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1766_
timestamp 0
transform 1 0 4416 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1767_
timestamp 0
transform 1 0 4968 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1768_
timestamp 0
transform 1 0 4876 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1769_
timestamp 0
transform 1 0 4324 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1770_
timestamp 0
transform 1 0 4140 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1771_
timestamp 0
transform -1 0 6072 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1772_
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 0
transform -1 0 4968 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1774_
timestamp 0
transform -1 0 3772 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1775__121
timestamp 0
transform -1 0 7452 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 0
transform 1 0 6808 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 0
transform -1 0 7544 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 0
transform -1 0 5612 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1778_
timestamp 0
transform -1 0 5704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1779_
timestamp 0
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1780_
timestamp 0
transform -1 0 4232 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1781_
timestamp 0
transform 1 0 4232 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1782_
timestamp 0
transform -1 0 5888 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1783_
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1784_
timestamp 0
transform 1 0 4508 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1785_
timestamp 0
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1786_
timestamp 0
transform 1 0 4784 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 0
transform 1 0 4600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1788_
timestamp 0
transform -1 0 5244 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1789__122
timestamp 0
transform -1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1790_
timestamp 0
transform -1 0 5428 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1791_
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1792_
timestamp 0
transform -1 0 9200 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1793_
timestamp 0
transform 1 0 6900 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1794_
timestamp 0
transform -1 0 6900 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1795_
timestamp 0
transform 1 0 6900 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1796_
timestamp 0
transform 1 0 8280 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1797_
timestamp 0
transform 1 0 7636 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1798_
timestamp 0
transform 1 0 7268 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1799_
timestamp 0
transform 1 0 7912 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1800_
timestamp 0
transform 1 0 7360 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 0
transform 1 0 8096 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 0
transform -1 0 7452 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1803__123
timestamp 0
transform -1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1803_
timestamp 0
transform 1 0 7452 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 0
transform -1 0 7452 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1805_
timestamp 0
transform 1 0 7360 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1806_
timestamp 0
transform -1 0 13248 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1807_
timestamp 0
transform -1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1808_
timestamp 0
transform -1 0 11960 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1809_
timestamp 0
transform -1 0 11868 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1810_
timestamp 0
transform -1 0 10672 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1811_
timestamp 0
transform -1 0 11316 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1812_
timestamp 0
transform -1 0 11408 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1813_
timestamp 0
transform 1 0 9292 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1814_
timestamp 0
transform 1 0 9752 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1815_
timestamp 0
transform 1 0 12144 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1816_
timestamp 0
transform 1 0 11960 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1817__124
timestamp 0
transform -1 0 10672 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 0
transform 1 0 9844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1818_
timestamp 0
transform 1 0 9568 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1820_
timestamp 0
transform -1 0 12144 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1821_
timestamp 0
transform 1 0 11868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1822_
timestamp 0
transform -1 0 11132 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1823_
timestamp 0
transform 1 0 10212 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1824_
timestamp 0
transform -1 0 9752 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1825_
timestamp 0
transform -1 0 10212 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1826_
timestamp 0
transform -1 0 10488 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1827_
timestamp 0
transform -1 0 9844 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1828_
timestamp 0
transform -1 0 11132 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1829_
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1830_
timestamp 0
transform 1 0 12328 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1831__125
timestamp 0
transform -1 0 10488 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1831_
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1832_
timestamp 0
transform 1 0 9384 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1833_
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  _1834_
timestamp 0
transform -1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _1835_
timestamp 0
transform -1 0 8004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _1836_
timestamp 0
transform 1 0 6532 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1837_
timestamp 0
transform 1 0 6992 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  _1838_
timestamp 0
transform -1 0 6532 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  _1839_
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1840_
timestamp 0
transform 1 0 6992 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  _1841_
timestamp 0
transform -1 0 8832 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1842_
timestamp 0
transform -1 0 8372 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1843_
timestamp 0
transform 1 0 6992 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1844_
timestamp 0
transform 1 0 6624 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1845__126
timestamp 0
transform -1 0 8740 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1845_
timestamp 0
transform 1 0 7636 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1846_
timestamp 0
transform 1 0 6808 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1847_
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1910_
timestamp 0
transform 1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1911_
timestamp 0
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1912_
timestamp 0
transform -1 0 8648 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1913_
timestamp 0
transform 1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1914_
timestamp 0
transform -1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1915_
timestamp 0
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1916_
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1917_
timestamp 0
transform 1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1918_
timestamp 0
transform -1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1919_
timestamp 0
transform 1 0 6992 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1920_
timestamp 0
transform 1 0 6072 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1921_
timestamp 0
transform 1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1922_
timestamp 0
transform 1 0 7176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1923_
timestamp 0
transform -1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1924_
timestamp 0
transform -1 0 9660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1925_
timestamp 0
transform -1 0 9936 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1926_
timestamp 0
transform -1 0 18124 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1927_
timestamp 0
transform -1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1928_
timestamp 0
transform -1 0 16100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1929_
timestamp 0
transform -1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1930_
timestamp 0
transform -1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1931_
timestamp 0
transform -1 0 19136 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1932_
timestamp 0
transform -1 0 18768 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1933_
timestamp 0
transform -1 0 14352 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1934_
timestamp 0
transform -1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1935_
timestamp 0
transform -1 0 17940 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1936_
timestamp 0
transform -1 0 18216 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1937_
timestamp 0
transform -1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1938_
timestamp 0
transform -1 0 17848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1939_
timestamp 0
transform -1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1940_
timestamp 0
transform -1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1941_
timestamp 0
transform -1 0 16928 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_23
timestamp 0
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_34
timestamp 0
transform 1 0 4232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_50
timestamp 0
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_62
timestamp 0
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_71
timestamp 0
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_76
timestamp 0
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_90
timestamp 0
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_104
timestamp 0
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_118
timestamp 0
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_132
timestamp 0
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 0
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_146
timestamp 0
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_162
timestamp 0
transform 1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 0
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_174
timestamp 0
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_188
timestamp 0
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 0
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_202
timestamp 0
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_216
timestamp 0
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 0
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_245
timestamp 0
transform 1 0 23644 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_35
timestamp 0
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52
timestamp 0
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_97
timestamp 0
transform 1 0 10028 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_101
timestamp 0
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 0
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_145
timestamp 0
transform 1 0 14444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 0
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_177
timestamp 0
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_195
timestamp 0
transform 1 0 19044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_207
timestamp 0
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_219
timestamp 0
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_237
timestamp 0
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 0
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_43
timestamp 0
transform 1 0 5060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_55
timestamp 0
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_67
timestamp 0
transform 1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_75
timestamp 0
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_93
timestamp 0
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_125
timestamp 0
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_137
timestamp 0
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_154
timestamp 0
transform 1 0 15272 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_166
timestamp 0
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_170
timestamp 0
transform 1 0 16744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_186
timestamp 0
transform 1 0 18216 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 0
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 0
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_233
timestamp 0
transform 1 0 22540 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_241
timestamp 0
transform 1 0 23276 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_50
timestamp 0
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 0
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_141
timestamp 0
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_163
timestamp 0
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_191
timestamp 0
transform 1 0 18676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_203
timestamp 0
transform 1 0 19780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_215
timestamp 0
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_237
timestamp 0
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_245
timestamp 0
transform 1 0 23644 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_37
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_55
timestamp 0
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_67
timestamp 0
transform 1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 0
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_112
timestamp 0
transform 1 0 11408 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_124
timestamp 0
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 0
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_149
timestamp 0
transform 1 0 14812 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_155
timestamp 0
transform 1 0 15364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_167
timestamp 0
transform 1 0 16468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_179
timestamp 0
transform 1 0 17572 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_191
timestamp 0
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 0
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_216
timestamp 0
transform 1 0 20976 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_228
timestamp 0
transform 1 0 22080 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_35
timestamp 0
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 0
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_73
timestamp 0
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_86
timestamp 0
transform 1 0 9016 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_98
timestamp 0
transform 1 0 10120 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_143
timestamp 0
transform 1 0 14260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_160
timestamp 0
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_187
timestamp 0
transform 1 0 18308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_199
timestamp 0
transform 1 0 19412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_203
timestamp 0
transform 1 0 19780 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 0
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_237
timestamp 0
transform 1 0 22908 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_37
timestamp 0
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_52
timestamp 0
transform 1 0 5888 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_64
timestamp 0
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_76
timestamp 0
transform 1 0 8096 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_101
timestamp 0
transform 1 0 10396 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_114
timestamp 0
transform 1 0 11592 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_129
timestamp 0
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_165
timestamp 0
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_173
timestamp 0
transform 1 0 17020 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_182
timestamp 0
transform 1 0 17848 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_190
timestamp 0
transform 1 0 18584 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_207
timestamp 0
transform 1 0 20148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_219
timestamp 0
transform 1 0 21252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_231
timestamp 0
transform 1 0 22356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_91
timestamp 0
transform 1 0 9476 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_121
timestamp 0
transform 1 0 12236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_146
timestamp 0
transform 1 0 14536 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_154
timestamp 0
transform 1 0 15272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_208
timestamp 0
transform 1 0 20240 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_220
timestamp 0
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_237
timestamp 0
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_35
timestamp 0
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_73
timestamp 0
transform 1 0 7820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 0
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 0
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_95
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_103
timestamp 0
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_125
timestamp 0
transform 1 0 12604 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 0
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_149
timestamp 0
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_160
timestamp 0
transform 1 0 15824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_164
timestamp 0
transform 1 0 16192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_186
timestamp 0
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_190
timestamp 0
transform 1 0 18584 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_209
timestamp 0
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_217
timestamp 0
transform 1 0 21068 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_230
timestamp 0
transform 1 0 22264 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_242
timestamp 0
transform 1 0 23368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_6
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_14
timestamp 0
transform 1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_29
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_47
timestamp 0
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 0
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_71
timestamp 0
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_76
timestamp 0
transform 1 0 8096 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_82
timestamp 0
transform 1 0 8648 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_91
timestamp 0
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_103
timestamp 0
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_142
timestamp 0
transform 1 0 14168 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_157
timestamp 0
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_164
timestamp 0
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_196
timestamp 0
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_208
timestamp 0
transform 1 0 20240 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_216
timestamp 0
transform 1 0 20976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_232
timestamp 0
transform 1 0 22448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_242
timestamp 0
transform 1 0 23368 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 0
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_54
timestamp 0
transform 1 0 6072 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_69
timestamp 0
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 0
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_103
timestamp 0
transform 1 0 10580 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_111
timestamp 0
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_123
timestamp 0
transform 1 0 12420 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_129
timestamp 0
transform 1 0 12972 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_150
timestamp 0
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_154
timestamp 0
transform 1 0 15272 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_160
timestamp 0
transform 1 0 15824 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_172
timestamp 0
transform 1 0 16928 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_184
timestamp 0
transform 1 0 18032 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_197
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_209
timestamp 0
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_245
timestamp 0
transform 1 0 23644 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_40
timestamp 0
transform 1 0 4784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_46
timestamp 0
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 0
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_120
timestamp 0
transform 1 0 12144 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_128
timestamp 0
transform 1 0 12880 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_140
timestamp 0
transform 1 0 13984 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_152
timestamp 0
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_156
timestamp 0
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_160
timestamp 0
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_172
timestamp 0
transform 1 0 16928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_180
timestamp 0
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_203
timestamp 0
transform 1 0 19780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_218
timestamp 0
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_235
timestamp 0
transform 1 0 22724 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_239
timestamp 0
transform 1 0 23092 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 0
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 0
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_71
timestamp 0
transform 1 0 7636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_113
timestamp 0
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_123
timestamp 0
transform 1 0 12420 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 0
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_168
timestamp 0
transform 1 0 16560 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_176
timestamp 0
transform 1 0 17296 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_182
timestamp 0
transform 1 0 17848 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 0
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 0
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 0
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_233
timestamp 0
transform 1 0 22540 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_241
timestamp 0
transform 1 0 23276 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_35
timestamp 0
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 0
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 0
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_72
timestamp 0
transform 1 0 7728 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_84
timestamp 0
transform 1 0 8832 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_97
timestamp 0
transform 1 0 10028 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 0
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_129
timestamp 0
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_142
timestamp 0
transform 1 0 14168 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_163
timestamp 0
transform 1 0 16100 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_172
timestamp 0
transform 1 0 16928 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_180
timestamp 0
transform 1 0 17664 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_186
timestamp 0
transform 1 0 18216 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_198
timestamp 0
transform 1 0 19320 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_210
timestamp 0
transform 1 0 20424 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 0
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_237
timestamp 0
transform 1 0 22908 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_6
timestamp 0
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_18
timestamp 0
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 0
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_59
timestamp 0
transform 1 0 6532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 0
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_164
timestamp 0
transform 1 0 16192 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_176
timestamp 0
transform 1 0 17296 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_183
timestamp 0
transform 1 0 17940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 0
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_220
timestamp 0
transform 1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_242
timestamp 0
transform 1 0 23368 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_6
timestamp 0
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_18
timestamp 0
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_30
timestamp 0
transform 1 0 3864 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_38
timestamp 0
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_52
timestamp 0
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_144
timestamp 0
transform 1 0 14352 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_152
timestamp 0
transform 1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_164
timestamp 0
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_193
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_201
timestamp 0
transform 1 0 19596 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_206
timestamp 0
transform 1 0 20056 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_216
timestamp 0
transform 1 0 20976 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_6
timestamp 0
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 0
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 0
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_44
timestamp 0
transform 1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_52
timestamp 0
transform 1 0 5888 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_64
timestamp 0
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_75
timestamp 0
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_91
timestamp 0
transform 1 0 9476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_101
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_127
timestamp 0
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_154
timestamp 0
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_172
timestamp 0
transform 1 0 16928 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_180
timestamp 0
transform 1 0 17664 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 0
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_209
timestamp 0
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_217
timestamp 0
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_229
timestamp 0
transform 1 0 22172 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_235
timestamp 0
transform 1 0 22724 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_239
timestamp 0
transform 1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_6
timestamp 0
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_18
timestamp 0
transform 1 0 2760 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_26
timestamp 0
transform 1 0 3496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 0
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_65
timestamp 0
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_79
timestamp 0
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_91
timestamp 0
transform 1 0 9476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_104
timestamp 0
transform 1 0 10672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_118
timestamp 0
transform 1 0 11960 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_132
timestamp 0
transform 1 0 13248 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_144
timestamp 0
transform 1 0 14352 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_152
timestamp 0
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_178
timestamp 0
transform 1 0 17480 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_184
timestamp 0
transform 1 0 18032 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_197
timestamp 0
transform 1 0 19228 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_208
timestamp 0
transform 1 0 20240 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_220
timestamp 0
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_237
timestamp 0
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_35
timestamp 0
transform 1 0 4324 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_45
timestamp 0
transform 1 0 5244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_57
timestamp 0
transform 1 0 6348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_104
timestamp 0
transform 1 0 10672 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_117
timestamp 0
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_125
timestamp 0
transform 1 0 12604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 0
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_157
timestamp 0
transform 1 0 15548 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_163
timestamp 0
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_168
timestamp 0
transform 1 0 16560 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_180
timestamp 0
transform 1 0 17664 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_192
timestamp 0
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_209
timestamp 0
transform 1 0 20332 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_219
timestamp 0
transform 1 0 21252 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_231
timestamp 0
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_243
timestamp 0
transform 1 0 23460 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_6
timestamp 0
transform 1 0 1656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_18
timestamp 0
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_30
timestamp 0
transform 1 0 3864 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_34
timestamp 0
transform 1 0 4232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_50
timestamp 0
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_88
timestamp 0
transform 1 0 9200 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_96
timestamp 0
transform 1 0 9936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_104
timestamp 0
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_133
timestamp 0
transform 1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_148
timestamp 0
transform 1 0 14720 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_160
timestamp 0
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_181
timestamp 0
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_189
timestamp 0
transform 1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_206
timestamp 0
transform 1 0 20056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 0
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_237
timestamp 0
transform 1 0 22908 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_6
timestamp 0
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_18
timestamp 0
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 0
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_61
timestamp 0
transform 1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_66
timestamp 0
transform 1 0 7176 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp 0
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_129
timestamp 0
transform 1 0 12972 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_149
timestamp 0
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_159
timestamp 0
transform 1 0 15732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_171
timestamp 0
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 0
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 0
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 0
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_202
timestamp 0
transform 1 0 19688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_217
timestamp 0
transform 1 0 21068 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_229
timestamp 0
transform 1 0 22172 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_241
timestamp 0
transform 1 0 23276 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_6
timestamp 0
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 0
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_30
timestamp 0
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_42
timestamp 0
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 0
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 0
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_120
timestamp 0
transform 1 0 12144 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_132
timestamp 0
transform 1 0 13248 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_150
timestamp 0
transform 1 0 14904 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_159
timestamp 0
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_185
timestamp 0
transform 1 0 18124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_197
timestamp 0
transform 1 0 19228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_209
timestamp 0
transform 1 0 20332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 0
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_237
timestamp 0
transform 1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_6
timestamp 0
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_18
timestamp 0
transform 1 0 2760 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_32
timestamp 0
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_46
timestamp 0
transform 1 0 5336 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_58
timestamp 0
transform 1 0 6440 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_75
timestamp 0
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_89
timestamp 0
transform 1 0 9292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_131
timestamp 0
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_150
timestamp 0
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_159
timestamp 0
transform 1 0 15732 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_171
timestamp 0
transform 1 0 16836 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_206
timestamp 0
transform 1 0 20056 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_218
timestamp 0
transform 1 0 21160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_231
timestamp 0
transform 1 0 22356 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_245
timestamp 0
transform 1 0 23644 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_40
timestamp 0
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp 0
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_63
timestamp 0
transform 1 0 6900 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_73
timestamp 0
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_85
timestamp 0
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 0
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_120
timestamp 0
transform 1 0 12144 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_132
timestamp 0
transform 1 0 13248 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_144
timestamp 0
transform 1 0 14352 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_156
timestamp 0
transform 1 0 15456 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_173
timestamp 0
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_179
timestamp 0
transform 1 0 17572 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_196
timestamp 0
transform 1 0 19136 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_208
timestamp 0
transform 1 0 20240 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_232
timestamp 0
transform 1 0 22448 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_245
timestamp 0
transform 1 0 23644 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_6
timestamp 0
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_18
timestamp 0
transform 1 0 2760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_22
timestamp 0
transform 1 0 3128 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_48
timestamp 0
transform 1 0 5520 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_71
timestamp 0
transform 1 0 7636 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_106
timestamp 0
transform 1 0 10856 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_118
timestamp 0
transform 1 0 11960 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_130
timestamp 0
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 0
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_162
timestamp 0
transform 1 0 16008 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_174
timestamp 0
transform 1 0 17112 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_180
timestamp 0
transform 1 0 17664 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_186
timestamp 0
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 0
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_209
timestamp 0
transform 1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_215
timestamp 0
transform 1 0 20884 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_230
timestamp 0
transform 1 0 22264 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_242
timestamp 0
transform 1 0 23368 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_6
timestamp 0
transform 1 0 1656 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_18
timestamp 0
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_30
timestamp 0
transform 1 0 3864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_36
timestamp 0
transform 1 0 4416 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_45
timestamp 0
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 0
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_63
timestamp 0
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_74
timestamp 0
transform 1 0 7912 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_86
timestamp 0
transform 1 0 9016 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_92
timestamp 0
transform 1 0 9568 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_102
timestamp 0
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 0
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_121
timestamp 0
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_131
timestamp 0
transform 1 0 13156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_139
timestamp 0
transform 1 0 13892 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_144
timestamp 0
transform 1 0 14352 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_156
timestamp 0
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_194
timestamp 0
transform 1 0 18952 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_206
timestamp 0
transform 1 0 20056 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_218
timestamp 0
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_232
timestamp 0
transform 1 0 22448 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_240
timestamp 0
transform 1 0 23184 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_6
timestamp 0
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_18
timestamp 0
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 0
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_37
timestamp 0
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_49
timestamp 0
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_61
timestamp 0
transform 1 0 6716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_74
timestamp 0
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 0
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_89
timestamp 0
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_102
timestamp 0
transform 1 0 10488 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_114
timestamp 0
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_135
timestamp 0
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_216
timestamp 0
transform 1 0 20976 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_228
timestamp 0
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_240
timestamp 0
transform 1 0 23184 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_6
timestamp 0
transform 1 0 1656 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_18
timestamp 0
transform 1 0 2760 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_30
timestamp 0
transform 1 0 3864 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_50
timestamp 0
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_63
timestamp 0
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_67
timestamp 0
transform 1 0 7268 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_79
timestamp 0
transform 1 0 8372 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_91
timestamp 0
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_103
timestamp 0
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_131
timestamp 0
transform 1 0 13156 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_143
timestamp 0
transform 1 0 14260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_151
timestamp 0
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_188
timestamp 0
transform 1 0 18400 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_192
timestamp 0
transform 1 0 18768 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_196
timestamp 0
transform 1 0 19136 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_208
timestamp 0
transform 1 0 20240 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_220
timestamp 0
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_237
timestamp 0
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_53
timestamp 0
transform 1 0 5980 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_89
timestamp 0
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_96
timestamp 0
transform 1 0 9936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_100
timestamp 0
transform 1 0 10304 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_110
timestamp 0
transform 1 0 11224 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_118
timestamp 0
transform 1 0 11960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_131
timestamp 0
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_147
timestamp 0
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_155
timestamp 0
transform 1 0 15364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_163
timestamp 0
transform 1 0 16100 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_173
timestamp 0
transform 1 0 17020 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_181
timestamp 0
transform 1 0 17756 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_185
timestamp 0
transform 1 0 18124 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 0
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_209
timestamp 0
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_217
timestamp 0
transform 1 0 21068 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_238
timestamp 0
transform 1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_242
timestamp 0
transform 1 0 23368 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_6
timestamp 0
transform 1 0 1656 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_18
timestamp 0
transform 1 0 2760 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_26
timestamp 0
transform 1 0 3496 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_43
timestamp 0
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_81
timestamp 0
transform 1 0 8556 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_92
timestamp 0
transform 1 0 9568 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_104
timestamp 0
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_120
timestamp 0
transform 1 0 12144 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_128
timestamp 0
transform 1 0 12880 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_135
timestamp 0
transform 1 0 13524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_141
timestamp 0
transform 1 0 14076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_164
timestamp 0
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_190
timestamp 0
transform 1 0 18584 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_198
timestamp 0
transform 1 0 19320 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 0
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_232
timestamp 0
transform 1 0 22448 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_245
timestamp 0
transform 1 0 23644 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_6
timestamp 0
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 0
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 0
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_46
timestamp 0
transform 1 0 5336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_54
timestamp 0
transform 1 0 6072 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_69
timestamp 0
transform 1 0 7452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 0
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_88
timestamp 0
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_93
timestamp 0
transform 1 0 9660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_105
timestamp 0
transform 1 0 10764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_134
timestamp 0
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_146
timestamp 0
transform 1 0 14536 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_152
timestamp 0
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_164
timestamp 0
transform 1 0 16192 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_176
timestamp 0
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_181
timestamp 0
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_188
timestamp 0
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_209
timestamp 0
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_217
timestamp 0
transform 1 0 21068 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_229
timestamp 0
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_245
timestamp 0
transform 1 0 23644 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_6
timestamp 0
transform 1 0 1656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_18
timestamp 0
transform 1 0 2760 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_26
timestamp 0
transform 1 0 3496 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_34
timestamp 0
transform 1 0 4232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_46
timestamp 0
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 0
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_81
timestamp 0
transform 1 0 8556 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_91
timestamp 0
transform 1 0 9476 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_103
timestamp 0
transform 1 0 10580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 0
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_181
timestamp 0
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_189
timestamp 0
transform 1 0 18492 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 0
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 0
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 0
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 0
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_237
timestamp 0
transform 1 0 22908 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 0
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_46
timestamp 0
transform 1 0 5336 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_54
timestamp 0
transform 1 0 6072 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_67
timestamp 0
transform 1 0 7268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_79
timestamp 0
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_107
timestamp 0
transform 1 0 10948 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_119
timestamp 0
transform 1 0 12052 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_131
timestamp 0
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_151
timestamp 0
transform 1 0 14996 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_159
timestamp 0
transform 1 0 15732 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_163
timestamp 0
transform 1 0 16100 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_174
timestamp 0
transform 1 0 17112 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_186
timestamp 0
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 0
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 0
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 0
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_233
timestamp 0
transform 1 0 22540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_241
timestamp 0
transform 1 0 23276 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_23
timestamp 0
transform 1 0 3220 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_40
timestamp 0
transform 1 0 4784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_52
timestamp 0
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_64
timestamp 0
transform 1 0 6992 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_76
timestamp 0
transform 1 0 8096 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_82
timestamp 0
transform 1 0 8648 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_95
timestamp 0
transform 1 0 9844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_106
timestamp 0
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_122
timestamp 0
transform 1 0 12328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_134
timestamp 0
transform 1 0 13432 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_159
timestamp 0
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_183
timestamp 0
transform 1 0 17940 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_191
timestamp 0
transform 1 0 18676 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_203
timestamp 0
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 0
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_237
timestamp 0
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_245
timestamp 0
transform 1 0 23644 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_6
timestamp 0
transform 1 0 1656 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_18
timestamp 0
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_26
timestamp 0
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_40
timestamp 0
transform 1 0 4784 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_48
timestamp 0
transform 1 0 5520 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_72
timestamp 0
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_92
timestamp 0
transform 1 0 9568 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_131
timestamp 0
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_147
timestamp 0
transform 1 0 14628 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 0
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_165
timestamp 0
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_169
timestamp 0
transform 1 0 16652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_182
timestamp 0
transform 1 0 17848 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_190
timestamp 0
transform 1 0 18584 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_222
timestamp 0
transform 1 0 21528 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_240
timestamp 0
transform 1 0 23184 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_6
timestamp 0
transform 1 0 1656 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_18
timestamp 0
transform 1 0 2760 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 0
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 0
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 0
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 0
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_81
timestamp 0
transform 1 0 8556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_90
timestamp 0
transform 1 0 9384 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_96
timestamp 0
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_108
timestamp 0
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_145
timestamp 0
transform 1 0 14444 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_151
timestamp 0
transform 1 0 14996 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 0
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_175
timestamp 0
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_187
timestamp 0
transform 1 0 18308 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_216
timestamp 0
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_237
timestamp 0
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_57
timestamp 0
transform 1 0 6348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_63
timestamp 0
transform 1 0 6900 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_75
timestamp 0
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 0
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_90
timestamp 0
transform 1 0 9384 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_102
timestamp 0
transform 1 0 10488 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_114
timestamp 0
transform 1 0 11592 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_118
timestamp 0
transform 1 0 11960 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_131
timestamp 0
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_158
timestamp 0
transform 1 0 15640 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_187
timestamp 0
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 0
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_233
timestamp 0
transform 1 0 22540 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_241
timestamp 0
transform 1 0 23276 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 0
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 0
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 0
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 0
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_70
timestamp 0
transform 1 0 7544 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_78
timestamp 0
transform 1 0 8280 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_100
timestamp 0
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_127
timestamp 0
transform 1 0 12788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_139
timestamp 0
transform 1 0 13892 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_153
timestamp 0
transform 1 0 15180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_165
timestamp 0
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_178
timestamp 0
transform 1 0 17480 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_190
timestamp 0
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_202
timestamp 0
transform 1 0 19688 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_218
timestamp 0
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_237
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 0
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_53
timestamp 0
transform 1 0 5980 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_69
timestamp 0
transform 1 0 7452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_81
timestamp 0
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_90
timestamp 0
transform 1 0 9384 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_102
timestamp 0
transform 1 0 10488 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_114
timestamp 0
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_126
timestamp 0
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 0
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_141
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_150
timestamp 0
transform 1 0 14904 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_162
timestamp 0
transform 1 0 16008 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_174
timestamp 0
transform 1 0 17112 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_186
timestamp 0
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 0
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 0
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 0
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 0
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_245
timestamp 0
transform 1 0 23644 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 0
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 0
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_75
timestamp 0
transform 1 0 8004 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_97
timestamp 0
transform 1 0 10028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_109
timestamp 0
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_137
timestamp 0
transform 1 0 13708 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 0
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 0
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_190
timestamp 0
transform 1 0 18584 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_202
timestamp 0
transform 1 0 19688 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_214
timestamp 0
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 0
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 0
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 0
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 0
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 0
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 0
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_88
timestamp 0
transform 1 0 9200 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_100
timestamp 0
transform 1 0 10304 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_112
timestamp 0
transform 1 0 11408 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_124
timestamp 0
transform 1 0 12512 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_136
timestamp 0
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_147
timestamp 0
transform 1 0 14628 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_151
timestamp 0
transform 1 0 14996 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_163
timestamp 0
transform 1 0 16100 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_175
timestamp 0
transform 1 0 17204 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_187
timestamp 0
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 0
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_221
timestamp 0
transform 1 0 21436 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_229
timestamp 0
transform 1 0 22172 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 0
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_27
timestamp 0
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_29
timestamp 0
transform 1 0 3772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_41
timestamp 0
transform 1 0 4876 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_49
timestamp 0
transform 1 0 5612 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 0
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_62
timestamp 0
transform 1 0 6808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_69
timestamp 0
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_76
timestamp 0
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_83
timestamp 0
transform 1 0 8740 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_85
timestamp 0
transform 1 0 8924 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_90
timestamp 0
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_97
timestamp 0
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_104
timestamp 0
transform 1 0 10672 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 0
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_118
timestamp 0
transform 1 0 11960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_125
timestamp 0
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_132
timestamp 0
transform 1 0 13248 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_139
timestamp 0
transform 1 0 13892 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_141
timestamp 0
transform 1 0 14076 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_146
timestamp 0
transform 1 0 14536 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_153
timestamp 0
transform 1 0 15180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_160
timestamp 0
transform 1 0 15824 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 0
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_174
timestamp 0
transform 1 0 17112 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_188
timestamp 0
transform 1 0 18400 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_197
timestamp 0
transform 1 0 19228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_209
timestamp 0
transform 1 0 20332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_216
timestamp 0
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_229
timestamp 0
transform 1 0 22172 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform -1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 6164 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform -1 0 8096 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform -1 0 12604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 12972 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform -1 0 23736 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 0
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 0
transform -1 0 18400 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 0
transform 1 0 23460 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 0
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 0
transform 1 0 23460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 0
transform 1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 0
transform 1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform -1 0 23736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 0
transform -1 0 23736 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 0
transform 1 0 23460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 0
transform 1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 0
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 0
transform 1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 0
transform 1 0 21344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 0
transform -1 0 6164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 0
transform 1 0 18768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 0
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 0
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 0
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 0
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 0
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input33
timestamp 0
transform -1 0 23736 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 0
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 0
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 0
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 0
transform -1 0 6808 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 0
transform -1 0 7452 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 0
transform -1 0 11960 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 0
transform -1 0 13892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 0
transform -1 0 23736 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 0
transform 1 0 14904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 0
transform -1 0 17756 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 0
transform -1 0 20976 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 0
transform -1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 0
transform 1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 0
transform 1 0 23460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 0
transform -1 0 23736 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 0
transform -1 0 23460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 0
transform -1 0 23736 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 0
transform 1 0 23460 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 0
transform 1 0 23460 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 0
transform 1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 0
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 0
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 0
transform -1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 0
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 0
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 0
transform -1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 0
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 0
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 0
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 0
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 0
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input66
timestamp 0
transform -1 0 23736 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 0
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input68
timestamp 0
transform -1 0 23736 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input69
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  output70
timestamp 0
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output71
timestamp 0
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output72
timestamp 0
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output73
timestamp 0
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output74
timestamp 0
transform -1 0 8740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output75
timestamp 0
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output76
timestamp 0
transform -1 0 9384 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output77
timestamp 0
transform -1 0 10672 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output78
timestamp 0
transform -1 0 10028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output79
timestamp 0
transform 1 0 23460 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output80
timestamp 0
transform -1 0 14536 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output81
timestamp 0
transform -1 0 16468 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output82
timestamp 0
transform 1 0 23460 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output83
timestamp 0
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output84
timestamp 0
transform 1 0 23184 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output85
timestamp 0
transform 1 0 23460 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output86
timestamp 0
transform 1 0 23460 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output87
timestamp 0
transform -1 0 15824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output88
timestamp 0
transform -1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output89
timestamp 0
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output90
timestamp 0
transform 1 0 23460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output91
timestamp 0
transform -1 0 20976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output92
timestamp 0
transform 1 0 23460 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output93
timestamp 0
transform -1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output94
timestamp 0
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output95
timestamp 0
transform -1 0 16468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output96
timestamp 0
transform 1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output97
timestamp 0
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output98
timestamp 0
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output99
timestamp 0
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output100
timestamp 0
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output101
timestamp 0
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output102
timestamp 0
transform -1 0 11316 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output103
timestamp 0
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output104
timestamp 0
transform -1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_42
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_43
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_44
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_45
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_46
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_47
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_48
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_49
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_50
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_51
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_52
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_53
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_54
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_55
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 24012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_56
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_57
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_58
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_59
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 24012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_60
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_61
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 24012 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_62
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_63
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 24012 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_64
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_65
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_66
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_67
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 24012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_68
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_69
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 24012 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_70
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_71
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 24012 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_72
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_73
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 0
transform -1 0 24012 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_74
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 0
transform -1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_75
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 0
transform -1 0 24012 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_76
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 0
transform -1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_77
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 0
transform -1 0 24012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_78
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 0
transform -1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_79
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 0
transform -1 0 24012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_80
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 0
transform -1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_81
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 0
transform -1 0 24012 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_82
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 0
transform -1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_83
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 0
transform -1 0 24012 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_90
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_91
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_94
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_95
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_108
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_109
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_110
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_112
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_113
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_114
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_115
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_117
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_118
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_119
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_123
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_136
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_137
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_138
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_142
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_143
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_146
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_147
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_150
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_151
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_153
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_154
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_155
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_157
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_158
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_159
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_162
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_163
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_167
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_188
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_190
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_191
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_192
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_194
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_195
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_196
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_197
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_199
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_201
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_202
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_203
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_204
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_205
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_206
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_207
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_208
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_209
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_210
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_211
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_214
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_215
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_216
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_217
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_218
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_219
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_220
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_221
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_222
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_223
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_224
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_230
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_231
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_233
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_234
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_235
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_236
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_237
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_238
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_239
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_242
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_243
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_244
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_245
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_246
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_247
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_248
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_249
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_250
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_251
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_252
timestamp 0
transform 1 0 3680 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_253
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_254
timestamp 0
transform 1 0 8832 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_255
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_256
timestamp 0
transform 1 0 13984 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_257
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_258
timestamp 0
transform 1 0 19136 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_259
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
<< labels >>
rlabel metal1 s 12558 25024 12558 25024 4 VGND
rlabel metal1 s 12558 24480 12558 24480 4 VPWR
rlabel metal1 s 14168 5746 14168 5746 4 _0030_
rlabel metal2 s 18216 14756 18216 14756 4 _0032_
rlabel metal1 s 17342 9656 17342 9656 4 _0033_
rlabel metal2 s 13294 9078 13294 9078 4 _0034_
rlabel metal2 s 13202 14348 13202 14348 4 _0035_
rlabel metal1 s 13800 10506 13800 10506 4 _0036_
rlabel metal1 s 14122 18598 14122 18598 4 _0037_
rlabel metal1 s 15640 8058 15640 8058 4 _0038_
rlabel metal1 s 8372 9418 8372 9418 4 _0039_
rlabel metal1 s 13570 10676 13570 10676 4 _0040_
rlabel metal1 s 14168 10778 14168 10778 4 _0041_
rlabel metal2 s 8050 9316 8050 9316 4 _0043_
rlabel metal2 s 6302 17476 6302 17476 4 _0044_
rlabel metal1 s 7038 18258 7038 18258 4 _0045_
rlabel metal2 s 7130 18224 7130 18224 4 _0046_
rlabel metal2 s 8970 18938 8970 18938 4 _0047_
rlabel metal2 s 9430 19210 9430 19210 4 _0048_
rlabel metal1 s 9706 17612 9706 17612 4 _0049_
rlabel metal2 s 17894 17850 17894 17850 4 _0050_
rlabel metal2 s 14122 20026 14122 20026 4 _0051_
rlabel metal2 s 15870 19380 15870 19380 4 _0052_
rlabel metal1 s 18446 19346 18446 19346 4 _0053_
rlabel metal1 s 9200 6766 9200 6766 4 _0054_
rlabel metal1 s 18170 18700 18170 18700 4 _0055_
rlabel metal1 s 19228 17170 19228 17170 4 _0056_
rlabel metal1 s 18400 16762 18400 16762 4 _0057_
rlabel metal2 s 14122 17374 14122 17374 4 _0058_
rlabel metal1 s 15640 8466 15640 8466 4 _0059_
rlabel metal2 s 17710 10506 17710 10506 4 _0060_
rlabel metal2 s 17986 9724 17986 9724 4 _0061_
rlabel metal2 s 16698 8262 16698 8262 4 _0062_
rlabel metal1 s 17526 8942 17526 8942 4 _0063_
rlabel metal1 s 15778 7378 15778 7378 4 _0064_
rlabel metal2 s 8418 6460 8418 6460 4 _0065_
rlabel metal1 s 15272 7378 15272 7378 4 _0066_
rlabel metal1 s 16698 9486 16698 9486 4 _0067_
rlabel metal1 s 7590 6766 7590 6766 4 _0068_
rlabel metal1 s 8418 7378 8418 7378 4 _0069_
rlabel metal1 s 5658 9520 5658 9520 4 _0070_
rlabel metal1 s 7544 9554 7544 9554 4 _0071_
rlabel metal1 s 9384 7378 9384 7378 4 _0072_
rlabel metal2 s 9430 17918 9430 17918 4 _0073_
rlabel metal1 s 6624 17782 6624 17782 4 _0074_
rlabel metal1 s 11109 8806 11109 8806 4 _0079_
rlabel metal1 s 10856 8602 10856 8602 4 _0080_
rlabel metal1 s 9476 8942 9476 8942 4 _0081_
rlabel metal1 s 10580 8806 10580 8806 4 _0082_
rlabel metal1 s 10442 8262 10442 8262 4 _0084_
rlabel metal1 s 9798 8806 9798 8806 4 _0085_
rlabel metal1 s 10212 8058 10212 8058 4 _0086_
rlabel metal1 s 10488 7990 10488 7990 4 _0087_
rlabel metal1 s 10672 5678 10672 5678 4 _0088_
rlabel metal1 s 11132 7922 11132 7922 4 _0090_
rlabel metal1 s 12052 8398 12052 8398 4 _0094_
rlabel metal1 s 8510 9044 8510 9044 4 _0105_
rlabel metal2 s 13386 7446 13386 7446 4 _0108_
rlabel metal1 s 8786 8874 8786 8874 4 _0111_
rlabel metal1 s 14329 7514 14329 7514 4 _0120_
rlabel metal2 s 12765 5882 12765 5882 4 _0121_
rlabel metal2 s 13938 8262 13938 8262 4 _0122_
rlabel metal1 s 13294 6766 13294 6766 4 _0123_
rlabel metal1 s 13110 7888 13110 7888 4 _0125_
rlabel metal1 s 13570 8058 13570 8058 4 _0126_
rlabel metal2 s 13478 6154 13478 6154 4 _0127_
rlabel metal1 s 13432 5610 13432 5610 4 _0128_
rlabel metal1 s 13432 6222 13432 6222 4 _0131_
rlabel metal1 s 13570 9146 13570 9146 4 _0146_
rlabel metal1 s 13340 8602 13340 8602 4 _0152_
rlabel metal1 s 4945 14246 4945 14246 4 _0161_
rlabel metal1 s 3519 14314 3519 14314 4 _0162_
rlabel metal1 s 4784 15130 4784 15130 4 _0163_
rlabel metal1 s 3634 14926 3634 14926 4 _0164_
rlabel metal1 s 3772 14994 3772 14994 4 _0166_
rlabel metal1 s 4370 15334 4370 15334 4 _0167_
rlabel metal2 s 3266 15878 3266 15878 4 _0168_
rlabel metal2 s 5106 15912 5106 15912 4 _0169_
rlabel metal1 s 3818 18292 3818 18292 4 _0170_
rlabel metal1 s 4508 16014 4508 16014 4 _0172_
rlabel metal2 s 5198 16218 5198 16218 4 _0176_
rlabel metal2 s 5474 15844 5474 15844 4 _0178_
rlabel metal1 s 4876 16762 4876 16762 4 _0187_
rlabel metal2 s 5014 16422 5014 16422 4 _0193_
rlabel metal2 s 4462 21148 4462 21148 4 _0202_
rlabel metal1 s 3703 21522 3703 21522 4 _0203_
rlabel metal2 s 4462 20026 4462 20026 4 _0204_
rlabel metal1 s 3680 20434 3680 20434 4 _0205_
rlabel metal2 s 4370 20842 4370 20842 4 _0207_
rlabel metal1 s 3910 19822 3910 19822 4 _0208_
rlabel metal1 s 4922 19856 4922 19856 4 _0209_
rlabel metal1 s 4646 18938 4646 18938 4 _0210_
rlabel metal1 s 5934 19822 5934 19822 4 _0211_
rlabel metal2 s 4002 18462 4002 18462 4 _0213_
rlabel metal1 s 4186 18224 4186 18224 4 _0217_
rlabel metal2 s 4278 18496 4278 18496 4 _0228_
rlabel metal1 s 4738 18734 4738 18734 4 _0234_
rlabel metal1 s 7061 22950 7061 22950 4 _0243_
rlabel metal1 s 7153 22746 7153 22746 4 _0244_
rlabel metal1 s 7130 20842 7130 20842 4 _0245_
rlabel metal1 s 6440 21454 6440 21454 4 _0246_
rlabel metal1 s 6302 21386 6302 21386 4 _0248_
rlabel metal1 s 6900 20978 6900 20978 4 _0249_
rlabel metal2 s 7314 21114 7314 21114 4 _0250_
rlabel metal1 s 7222 20570 7222 20570 4 _0251_
rlabel metal1 s 8418 20910 8418 20910 4 _0252_
rlabel metal1 s 6578 20434 6578 20434 4 _0254_
rlabel metal1 s 6992 19482 6992 19482 4 _0258_
rlabel metal2 s 6670 18972 6670 18972 4 _0269_
rlabel metal2 s 6762 19754 6762 19754 4 _0275_
rlabel metal1 s 9637 23698 9637 23698 4 _0284_
rlabel metal2 s 8418 23936 8418 23936 4 _0285_
rlabel metal1 s 9384 22202 9384 22202 4 _0286_
rlabel metal1 s 9108 23086 9108 23086 4 _0287_
rlabel metal1 s 8924 23086 8924 23086 4 _0289_
rlabel metal2 s 9522 22848 9522 22848 4 _0290_
rlabel metal1 s 10120 22406 10120 22406 4 _0291_
rlabel metal1 s 9522 21522 9522 21522 4 _0292_
rlabel metal1 s 12742 21080 12742 21080 4 _0293_
rlabel metal1 s 9062 21522 9062 21522 4 _0295_
rlabel metal1 s 9338 20570 9338 20570 4 _0299_
rlabel metal2 s 8970 19856 8970 19856 4 _0310_
rlabel metal2 s 9062 20944 9062 20944 4 _0316_
rlabel metal1 s 12765 21862 12765 21862 4 _0325_
rlabel metal1 s 12397 22610 12397 22610 4 _0326_
rlabel metal2 s 11822 21114 11822 21114 4 _0327_
rlabel metal1 s 12466 20876 12466 20876 4 _0328_
rlabel metal1 s 11868 22406 11868 22406 4 _0330_
rlabel metal2 s 11914 21148 11914 21148 4 _0331_
rlabel metal2 s 12650 20638 12650 20638 4 _0332_
rlabel metal2 s 13110 20604 13110 20604 4 _0333_
rlabel metal2 s 12742 19482 12742 19482 4 _0334_
rlabel metal1 s 12673 20978 12673 20978 4 _0336_
rlabel metal1 s 10626 19754 10626 19754 4 _0340_
rlabel metal1 s 9982 19686 9982 19686 4 _0351_
rlabel metal1 s 10580 19822 10580 19822 4 _0357_
rlabel metal1 s 13133 16422 13133 16422 4 _0366_
rlabel metal1 s 12880 16218 12880 16218 4 _0367_
rlabel metal1 s 12236 17170 12236 17170 4 _0368_
rlabel metal2 s 12650 17408 12650 17408 4 _0369_
rlabel metal2 s 12374 16388 12374 16388 4 _0371_
rlabel metal1 s 12052 16762 12052 16762 4 _0372_
rlabel metal2 s 13110 18054 13110 18054 4 _0373_
rlabel metal2 s 13294 18462 13294 18462 4 _0374_
rlabel metal1 s 13846 18122 13846 18122 4 _0375_
rlabel metal2 s 12650 18326 12650 18326 4 _0377_
rlabel metal1 s 12144 18734 12144 18734 4 _0381_
rlabel metal1 s 11224 17646 11224 17646 4 _0392_
rlabel metal1 s 11224 17306 11224 17306 4 _0398_
rlabel metal2 s 15962 16796 15962 16796 4 _0407_
rlabel metal1 s 15801 17170 15801 17170 4 _0408_
rlabel metal1 s 16330 17578 16330 17578 4 _0409_
rlabel metal2 s 15870 17204 15870 17204 4 _0410_
rlabel metal1 s 15180 17646 15180 17646 4 _0412_
rlabel metal1 s 16560 17714 16560 17714 4 _0413_
rlabel metal2 s 15318 18530 15318 18530 4 _0414_
rlabel metal2 s 14582 18530 14582 18530 4 _0415_
rlabel metal1 s 14674 19822 14674 19822 4 _0416_
rlabel metal1 s 14582 18190 14582 18190 4 _0418_
rlabel metal1 s 15226 18258 15226 18258 4 _0422_
rlabel metal1 s 17526 18394 17526 18394 4 _0433_
rlabel metal1 s 17158 17850 17158 17850 4 _0439_
rlabel metal2 s 15594 23936 15594 23936 4 _0448_
rlabel metal2 s 14743 23290 14743 23290 4 _0449_
rlabel metal1 s 14628 21998 14628 21998 4 _0450_
rlabel metal1 s 14996 22678 14996 22678 4 _0451_
rlabel metal2 s 14306 23018 14306 23018 4 _0453_
rlabel metal1 s 14720 21862 14720 21862 4 _0454_
rlabel metal1 s 15134 21522 15134 21522 4 _0455_
rlabel metal2 s 15134 21284 15134 21284 4 _0456_
rlabel metal2 s 16974 21114 16974 21114 4 _0457_
rlabel metal1 s 14812 20910 14812 20910 4 _0459_
rlabel metal2 s 14950 20230 14950 20230 4 _0463_
rlabel metal1 s 14674 20332 14674 20332 4 _0474_
rlabel metal2 s 14214 21216 14214 21216 4 _0480_
rlabel metal1 s 17986 23086 17986 23086 4 _0489_
rlabel metal1 s 17917 23698 17917 23698 4 _0490_
rlabel metal1 s 17342 22406 17342 22406 4 _0491_
rlabel metal1 s 17342 22610 17342 22610 4 _0492_
rlabel metal2 s 17066 23018 17066 23018 4 _0494_
rlabel metal1 s 16560 21930 16560 21930 4 _0495_
rlabel metal1 s 17802 21522 17802 21522 4 _0496_
rlabel metal1 s 17940 21114 17940 21114 4 _0497_
rlabel metal1 s 18952 21522 18952 21522 4 _0498_
rlabel metal2 s 17618 21522 17618 21522 4 _0500_
rlabel metal1 s 17296 20570 17296 20570 4 _0504_
rlabel metal2 s 16790 20060 16790 20060 4 _0515_
rlabel metal2 s 16698 20842 16698 20842 4 _0521_
rlabel metal1 s 22793 20774 22793 20774 4 _0530_
rlabel metal1 s 20769 22610 20769 22610 4 _0531_
rlabel metal1 s 21068 20842 21068 20842 4 _0532_
rlabel metal1 s 21206 20400 21206 20400 4 _0533_
rlabel metal1 s 20516 22406 20516 22406 4 _0535_
rlabel metal1 s 20884 20570 20884 20570 4 _0536_
rlabel metal2 s 20562 20910 20562 20910 4 _0537_
rlabel metal1 s 20792 20434 20792 20434 4 _0538_
rlabel metal1 s 20838 18258 20838 18258 4 _0539_
rlabel metal1 s 19826 21454 19826 21454 4 _0541_
rlabel metal2 s 19826 21114 19826 21114 4 _0545_
rlabel metal2 s 19458 20672 19458 20672 4 _0556_
rlabel metal1 s 19458 20502 19458 20502 4 _0562_
rlabel metal1 s 12213 3366 12213 3366 4 _0571_
rlabel metal1 s 10189 3162 10189 3162 4 _0572_
rlabel metal2 s 10718 3910 10718 3910 4 _0573_
rlabel metal1 s 11224 3570 11224 3570 4 _0574_
rlabel metal1 s 10764 4590 10764 4590 4 _0576_
rlabel metal1 s 10350 4046 10350 4046 4 _0577_
rlabel metal2 s 11362 4998 11362 4998 4 _0578_
rlabel metal1 s 11040 5270 11040 5270 4 _0579_
rlabel metal1 s 9660 5066 9660 5066 4 _0580_
rlabel metal1 s 10856 5746 10856 5746 4 _0582_
rlabel metal1 s 10994 5882 10994 5882 4 _0586_
rlabel metal1 s 10350 6426 10350 6426 4 _0597_
rlabel metal1 s 10212 3978 10212 3978 4 _0603_
rlabel metal1 s 23253 18258 23253 18258 4 _0612_
rlabel metal1 s 23253 18598 23253 18598 4 _0613_
rlabel metal2 s 22126 18258 22126 18258 4 _0614_
rlabel metal1 s 22126 18156 22126 18156 4 _0615_
rlabel metal1 s 22402 18258 22402 18258 4 _0617_
rlabel metal1 s 22678 17850 22678 17850 4 _0618_
rlabel metal1 s 21620 17578 21620 17578 4 _0619_
rlabel metal2 s 21390 17850 21390 17850 4 _0620_
rlabel metal2 s 22218 15844 22218 15844 4 _0621_
rlabel metal1 s 21528 18190 21528 18190 4 _0623_
rlabel metal1 s 20378 18224 20378 18224 4 _0627_
rlabel metal2 s 19550 18496 19550 18496 4 _0638_
rlabel metal1 s 20516 18666 20516 18666 4 _0644_
rlabel metal1 s 23253 14246 23253 14246 4 _0653_
rlabel metal1 s 23253 14994 23253 14994 4 _0654_
rlabel metal1 s 21114 15130 21114 15130 4 _0655_
rlabel metal1 s 22126 14994 22126 14994 4 _0656_
rlabel metal1 s 22218 14892 22218 14892 4 _0658_
rlabel metal2 s 21482 14960 21482 14960 4 _0659_
rlabel metal1 s 21804 14586 21804 14586 4 _0660_
rlabel metal1 s 21528 15062 21528 15062 4 _0661_
rlabel metal1 s 20102 14994 20102 14994 4 _0662_
rlabel metal2 s 22034 15198 22034 15198 4 _0664_
rlabel metal1 s 21850 16048 21850 16048 4 _0668_
rlabel metal1 s 20194 16218 20194 16218 4 _0679_
rlabel metal1 s 20470 15674 20470 15674 4 _0685_
rlabel metal1 s 19389 14314 19389 14314 4 _0694_
rlabel metal2 s 17181 13498 17181 13498 4 _0695_
rlabel metal2 s 18078 14518 18078 14518 4 _0696_
rlabel metal1 s 18262 14280 18262 14280 4 _0697_
rlabel metal2 s 17618 14620 17618 14620 4 _0699_
rlabel metal2 s 18446 14756 18446 14756 4 _0700_
rlabel metal2 s 17342 14586 17342 14586 4 _0701_
rlabel metal2 s 17158 14858 17158 14858 4 _0702_
rlabel metal1 s 16238 14382 16238 14382 4 _0703_
rlabel metal2 s 17986 15028 17986 15028 4 _0705_
rlabel metal2 s 18538 15504 18538 15504 4 _0709_
rlabel metal1 s 18078 16218 18078 16218 4 _0720_
rlabel metal1 s 18262 15130 18262 15130 4 _0726_
rlabel metal1 s 14237 12750 14237 12750 4 _0735_
rlabel metal1 s 13777 13226 13777 13226 4 _0736_
rlabel metal1 s 14352 14042 14352 14042 4 _0737_
rlabel metal1 s 14076 13838 14076 13838 4 _0738_
rlabel metal2 s 13846 14110 13846 14110 4 _0740_
rlabel metal1 s 14168 14246 14168 14246 4 _0741_
rlabel metal1 s 15042 13226 15042 13226 4 _0742_
rlabel metal1 s 15640 13294 15640 13294 4 _0743_
rlabel metal1 s 15778 13158 15778 13158 4 _0744_
rlabel metal1 s 15548 13906 15548 13906 4 _0746_
rlabel metal2 s 15134 14671 15134 14671 4 _0750_
rlabel metal1 s 14766 15334 14766 15334 4 _0761_
rlabel metal1 s 14674 14586 14674 14586 4 _0767_
rlabel metal2 s 17158 11968 17158 11968 4 _0776_
rlabel metal1 s 14789 11050 14789 11050 4 _0777_
rlabel metal1 s 15962 10030 15962 10030 4 _0778_
rlabel metal1 s 15686 11696 15686 11696 4 _0779_
rlabel metal2 s 15594 12002 15594 12002 4 _0781_
rlabel metal2 s 15870 10268 15870 10268 4 _0782_
rlabel metal2 s 16514 11662 16514 11662 4 _0783_
rlabel metal1 s 16560 11118 16560 11118 4 _0784_
rlabel metal2 s 18538 11526 18538 11526 4 _0785_
rlabel metal2 s 15962 11356 15962 11356 4 _0787_
rlabel metal1 s 16238 8874 16238 8874 4 _0791_
rlabel metal2 s 15778 9316 15778 9316 4 _0802_
rlabel metal1 s 15548 9690 15548 9690 4 _0808_
rlabel metal1 s 21045 12614 21045 12614 4 _0817_
rlabel metal2 s 20746 13056 20746 13056 4 _0818_
rlabel metal2 s 19182 13056 19182 13056 4 _0819_
rlabel metal1 s 19642 12886 19642 12886 4 _0820_
rlabel metal2 s 20010 13124 20010 13124 4 _0822_
rlabel metal1 s 19458 12818 19458 12818 4 _0823_
rlabel metal2 s 20194 11934 20194 11934 4 _0824_
rlabel metal1 s 19596 11730 19596 11730 4 _0825_
rlabel metal2 s 20746 11084 20746 11084 4 _0826_
rlabel metal2 s 18998 12002 18998 12002 4 _0828_
rlabel metal2 s 18446 11152 18446 11152 4 _0832_
rlabel metal1 s 18216 10778 18216 10778 4 _0843_
rlabel metal1 s 18538 12614 18538 12614 4 _0849_
rlabel metal2 s 23046 10540 23046 10540 4 _0858_
rlabel metal1 s 23345 10642 23345 10642 4 _0859_
rlabel metal2 s 22126 10438 22126 10438 4 _0860_
rlabel metal1 s 22448 10030 22448 10030 4 _0861_
rlabel metal2 s 22678 10268 22678 10268 4 _0863_
rlabel metal2 s 22034 10404 22034 10404 4 _0864_
rlabel metal1 s 21712 11050 21712 11050 4 _0865_
rlabel metal1 s 21390 10234 21390 10234 4 _0866_
rlabel metal1 s 22126 7956 22126 7956 4 _0867_
rlabel metal1 s 20976 10574 20976 10574 4 _0869_
rlabel metal2 s 20470 10234 20470 10234 4 _0873_
rlabel metal1 s 19918 9894 19918 9894 4 _0884_
rlabel metal2 s 19642 10268 19642 10268 4 _0890_
rlabel metal1 s 23253 7718 23253 7718 4 _0899_
rlabel metal2 s 23046 7888 23046 7888 4 _0900_
rlabel metal2 s 22218 8058 22218 8058 4 _0901_
rlabel metal1 s 22356 8058 22356 8058 4 _0902_
rlabel metal1 s 22678 8432 22678 8432 4 _0904_
rlabel metal2 s 21758 8092 21758 8092 4 _0905_
rlabel metal1 s 21804 6698 21804 6698 4 _0906_
rlabel metal2 s 22494 7242 22494 7242 4 _0907_
rlabel metal1 s 20240 6834 20240 6834 4 _0908_
rlabel metal1 s 22310 7820 22310 7820 4 _0910_
rlabel metal2 s 21114 7514 21114 7514 4 _0914_
rlabel metal1 s 20240 7718 20240 7718 4 _0925_
rlabel metal1 s 20608 7786 20608 7786 4 _0931_
rlabel metal2 s 20907 4794 20907 4794 4 _0940_
rlabel metal1 s 20447 4794 20447 4794 4 _0941_
rlabel metal1 s 18952 5882 18952 5882 4 _0942_
rlabel metal1 s 20056 5610 20056 5610 4 _0943_
rlabel metal1 s 20056 5678 20056 5678 4 _0945_
rlabel metal1 s 19504 5882 19504 5882 4 _0946_
rlabel metal1 s 19274 5780 19274 5780 4 _0947_
rlabel metal2 s 18538 6494 18538 6494 4 _0948_
rlabel metal2 s 17618 5882 17618 5882 4 _0949_
rlabel metal2 s 18906 6460 18906 6460 4 _0951_
rlabel metal2 s 19090 7888 19090 7888 4 _0955_
rlabel metal1 s 18538 8602 18538 8602 4 _0966_
rlabel metal1 s 18538 6426 18538 6426 4 _0972_
rlabel metal2 s 18837 3162 18837 3162 4 _0981_
rlabel metal1 s 18377 3026 18377 3026 4 _0982_
rlabel metal1 s 17250 3706 17250 3706 4 _0983_
rlabel metal2 s 18354 3876 18354 3876 4 _0984_
rlabel metal2 s 18170 3774 18170 3774 4 _0986_
rlabel metal1 s 17756 3706 17756 3706 4 _0987_
rlabel metal1 s 17802 3570 17802 3570 4 _0988_
rlabel metal1 s 17940 5270 17940 5270 4 _0989_
rlabel metal1 s 15410 5134 15410 5134 4 _0990_
rlabel metal1 s 17848 5134 17848 5134 4 _0992_
rlabel metal2 s 17250 6256 17250 6256 4 _0996_
rlabel metal1 s 16974 6630 16974 6630 4 _1007_
rlabel metal1 s 16974 3978 16974 3978 4 _1013_
rlabel metal1 s 8165 3026 8165 3026 4 _1022_
rlabel metal1 s 7291 2618 7291 2618 4 _1023_
rlabel metal2 s 8142 4352 8142 4352 4 _1024_
rlabel metal1 s 7498 4046 7498 4046 4 _1025_
rlabel metal1 s 6670 4080 6670 4080 4 _1027_
rlabel metal2 s 7958 3876 7958 3876 4 _1028_
rlabel metal1 s 7268 4250 7268 4250 4 _1029_
rlabel metal1 s 7866 4590 7866 4590 4 _1030_
rlabel metal1 s 5934 4624 5934 4624 4 _1031_
rlabel metal1 s 7866 5134 7866 5134 4 _1033_
rlabel metal1 s 8418 5134 8418 5134 4 _1037_
rlabel metal1 s 8418 6426 8418 6426 4 _1048_
rlabel metal2 s 8510 5134 8510 5134 4 _1054_
rlabel metal1 s 15663 2618 15663 2618 4 _1063_
rlabel metal1 s 15065 2618 15065 2618 4 _1064_
rlabel metal1 s 15640 4114 15640 4114 4 _1065_
rlabel metal1 s 15686 3162 15686 3162 4 _1066_
rlabel metal2 s 14858 3672 14858 3672 4 _1068_
rlabel metal2 s 15226 3723 15226 3723 4 _1069_
rlabel metal2 s 14766 4454 14766 4454 4 _1070_
rlabel metal1 s 14766 4794 14766 4794 4 _1071_
rlabel metal1 s 14996 4590 14996 4590 4 _1074_
rlabel metal2 s 15778 5712 15778 5712 4 _1078_
rlabel metal1 s 15456 6426 15456 6426 4 _1089_
rlabel metal2 s 15594 3995 15594 3995 4 _1095_
rlabel metal1 s 5497 3026 5497 3026 4 _1104_
rlabel metal1 s 4922 2482 4922 2482 4 _1105_
rlabel metal1 s 3956 4114 3956 4114 4 _1106_
rlabel metal2 s 4830 3298 4830 3298 4 _1107_
rlabel metal1 s 4784 3502 4784 3502 4 _1109_
rlabel metal2 s 5014 4080 5014 4080 4 _1110_
rlabel metal1 s 4462 4250 4462 4250 4 _1111_
rlabel metal1 s 5060 4250 5060 4250 4 _1112_
rlabel metal1 s 5198 5270 5198 5270 4 _1113_
rlabel metal1 s 5658 4114 5658 4114 4 _1115_
rlabel metal1 s 5520 4794 5520 4794 4 _1119_
rlabel metal2 s 5106 5440 5106 5440 4 _1130_
rlabel metal1 s 5336 4454 5336 4454 4 _1136_
rlabel metal1 s 4255 7378 4255 7378 4 _1145_
rlabel metal1 s 3059 7378 3059 7378 4 _1146_
rlabel metal1 s 5014 6970 5014 6970 4 _1147_
rlabel metal1 s 4738 6834 4738 6834 4 _1148_
rlabel metal2 s 4370 7684 4370 7684 4 _1150_
rlabel metal1 s 5244 7514 5244 7514 4 _1151_
rlabel metal1 s 4830 8466 4830 8466 4 _1152_
rlabel metal2 s 5658 8262 5658 8262 4 _1153_
rlabel metal2 s 5474 9554 5474 9554 4 _1154_
rlabel metal1 s 5290 7854 5290 7854 4 _1156_
rlabel metal1 s 6210 7344 6210 7344 4 _1160_
rlabel metal1 s 6946 7174 6946 7174 4 _1171_
rlabel metal1 s 5566 7752 5566 7752 4 _1177_
rlabel metal1 s 5313 12818 5313 12818 4 _1186_
rlabel metal1 s 4623 12682 4623 12682 4 _1187_
rlabel metal1 s 4462 11798 4462 11798 4 _1188_
rlabel metal1 s 4416 11730 4416 11730 4 _1189_
rlabel metal2 s 5566 11866 5566 11866 4 _1191_
rlabel metal1 s 4922 11662 4922 11662 4 _1192_
rlabel metal2 s 5842 11322 5842 11322 4 _1193_
rlabel metal1 s 5750 10778 5750 10778 4 _1194_
rlabel metal1 s 6187 11186 6187 11186 4 _1195_
rlabel metal2 s 5106 10880 5106 10880 4 _1197_
rlabel metal2 s 5290 10234 5290 10234 4 _1201_
rlabel metal2 s 4922 9792 4922 9792 4 _1212_
rlabel metal2 s 5014 10574 5014 10574 4 _1218_
rlabel metal1 s 8809 12818 8809 12818 4 _1227_
rlabel metal2 s 6946 13056 6946 13056 4 _1228_
rlabel metal1 s 7222 12104 7222 12104 4 _1229_
rlabel metal1 s 6670 12172 6670 12172 4 _1230_
rlabel metal1 s 6946 12274 6946 12274 4 _1232_
rlabel metal1 s 7590 12206 7590 12206 4 _1233_
rlabel metal1 s 8188 12682 8188 12682 4 _1234_
rlabel metal1 s 8418 11866 8418 11866 4 _1235_
rlabel metal1 s 9016 12274 9016 12274 4 _1236_
rlabel metal1 s 7774 11526 7774 11526 4 _1238_
rlabel metal2 s 7866 10608 7866 10608 4 _1242_
rlabel metal1 s 7222 9962 7222 9962 4 _1253_
rlabel metal1 s 7222 10030 7222 10030 4 _1259_
rlabel metal1 s 12857 11730 12857 11730 4 _1268_
rlabel metal2 s 12466 11628 12466 11628 4 _1269_
rlabel metal2 s 11546 11322 11546 11322 4 _1270_
rlabel metal1 s 11960 11662 11960 11662 4 _1271_
rlabel metal2 s 11914 11458 11914 11458 4 _1273_
rlabel metal1 s 11546 11186 11546 11186 4 _1274_
rlabel metal1 s 10764 12818 10764 12818 4 _1275_
rlabel metal1 s 10074 12410 10074 12410 4 _1276_
rlabel metal1 s 9890 14450 9890 14450 4 _1277_
rlabel metal1 s 10074 12308 10074 12308 4 _1279_
rlabel metal1 s 10166 11866 10166 11866 4 _1283_
rlabel metal2 s 10074 11356 10074 11356 4 _1294_
rlabel metal1 s 9982 11186 9982 11186 4 _1300_
rlabel metal2 s 11983 14042 11983 14042 4 _1309_
rlabel metal2 s 12834 14620 12834 14620 4 _1310_
rlabel metal2 s 10718 15266 10718 15266 4 _1311_
rlabel metal2 s 10902 14756 10902 14756 4 _1312_
rlabel metal1 s 11730 14858 11730 14858 4 _1314_
rlabel metal2 s 10626 15232 10626 15232 4 _1315_
rlabel metal1 s 9752 14994 9752 14994 4 _1316_
rlabel metal2 s 9430 14790 9430 14790 4 _1317_
rlabel metal2 s 8786 15334 8786 15334 4 _1318_
rlabel metal1 s 10350 14518 10350 14518 4 _1320_
rlabel metal1 s 10304 14586 10304 14586 4 _1324_
rlabel metal1 s 9798 16218 9798 16218 4 _1335_
rlabel metal1 s 9982 15674 9982 15674 4 _1341_
rlabel metal2 s 7521 14586 7521 14586 4 _1350_
rlabel metal1 s 7475 14246 7475 14246 4 _1351_
rlabel metal2 s 6946 16048 6946 16048 4 _1352_
rlabel metal1 s 7452 16082 7452 16082 4 _1353_
rlabel metal1 s 6624 15538 6624 15538 4 _1355_
rlabel metal1 s 7498 16218 7498 16218 4 _1356_
rlabel metal2 s 6486 15640 6486 15640 4 _1357_
rlabel metal1 s 6486 15470 6486 15470 4 _1358_
rlabel metal1 s 7820 15538 7820 15538 4 _1361_
rlabel metal1 s 7912 15674 7912 15674 4 _1365_
rlabel metal1 s 7498 17510 7498 17510 4 _1376_
rlabel metal1 s 7176 16762 7176 16762 4 _1382_
rlabel metal2 s 3266 1588 3266 1588 4 a[0]
rlabel metal3 s 1050 13668 1050 13668 4 a[10]
rlabel metal3 s 1050 20468 1050 20468 4 a[11]
rlabel metal1 s 5888 24786 5888 24786 4 a[12]
rlabel metal1 s 7820 24786 7820 24786 4 a[13]
rlabel metal1 s 12328 24786 12328 24786 4 a[14]
rlabel metal1 s 12972 24786 12972 24786 4 a[15]
rlabel metal1 s 23552 23698 23552 23698 4 a[16]
rlabel metal1 s 16928 24786 16928 24786 4 a[17]
rlabel metal1 s 18124 24786 18124 24786 4 a[18]
rlabel metal2 s 23690 22559 23690 22559 4 a[19]
rlabel metal2 s 11638 1588 11638 1588 4 a[1]
rlabel metal2 s 23690 21913 23690 21913 4 a[20]
rlabel metal2 s 23690 16473 23690 16473 4 a[21]
rlabel metal1 s 23552 15470 23552 15470 4 a[22]
rlabel metal2 s 23690 5015 23690 5015 4 a[23]
rlabel metal2 s 23690 11679 23690 11679 4 a[24]
rlabel metal1 s 23552 12818 23552 12818 4 a[25]
rlabel metal1 s 23552 5678 23552 5678 4 a[26]
rlabel metal2 s 23690 6239 23690 6239 4 a[27]
rlabel metal2 s 23690 2907 23690 2907 4 a[28]
rlabel metal2 s 21298 1588 21298 1588 4 a[29]
rlabel metal2 s 5842 1588 5842 1588 4 a[2]
rlabel metal2 s 18722 1588 18722 1588 4 a[30]
rlabel metal2 s 14858 1554 14858 1554 4 a[31]
rlabel metal2 s 3910 1588 3910 1588 4 a[3]
rlabel metal3 s 1050 6868 1050 6868 4 a[4]
rlabel metal3 s 1050 10948 1050 10948 4 a[5]
rlabel metal3 s 0 12928 800 13048 4 a[6]
port 31 nsew
rlabel metal2 s 12926 1588 12926 1588 4 a[7]
rlabel metal3 s 0 17008 800 17128 4 a[8]
port 33 nsew
rlabel metal3 s 0 15648 800 15768 4 a[9]
port 34 nsew
rlabel metal2 s 23690 24667 23690 24667 4 ainv
rlabel metal2 s 10350 823 10350 823 4 b[0]
rlabel metal3 s 0 14288 800 14408 4 b[10]
port 37 nsew
rlabel metal3 s 0 21088 800 21208 4 b[11]
port 38 nsew
rlabel metal1 s 6532 24786 6532 24786 4 b[12]
rlabel metal1 s 7176 24786 7176 24786 4 b[13]
rlabel metal1 s 11684 24786 11684 24786 4 b[14]
rlabel metal1 s 13708 24786 13708 24786 4 b[15]
rlabel metal1 s 23506 19346 23506 19346 4 b[16]
rlabel metal1 s 14996 24786 14996 24786 4 b[17]
rlabel metal1 s 17480 24786 17480 24786 4 b[18]
rlabel metal1 s 20700 24786 20700 24786 4 b[19]
rlabel metal2 s 5198 1554 5198 1554 4 b[1]
rlabel metal1 s 23552 20910 23552 20910 4 b[20]
rlabel metal2 s 23690 15895 23690 15895 4 b[21]
rlabel metal2 s 23690 14127 23690 14127 4 b[22]
rlabel metal2 s 23414 13787 23414 13787 4 b[23]
rlabel metal1 s 23552 11118 23552 11118 4 b[24]
rlabel metal2 s 23690 13141 23690 13141 4 b[25]
rlabel metal2 s 23690 10149 23690 10149 4 b[26]
rlabel metal2 s 23690 7463 23690 7463 4 b[27]
rlabel metal3 s 23690 3485 23690 3485 4 b[28]
rlabel metal2 s 19366 1588 19366 1588 4 b[29]
rlabel metal2 s 7130 1588 7130 1588 4 b[2]
rlabel metal2 s 17434 1588 17434 1588 4 b[30]
rlabel metal2 s 14214 1588 14214 1588 4 b[31]
rlabel metal2 s 4554 1027 4554 1027 4 b[3]
rlabel metal3 s 0 7488 800 7608 4 b[4]
port 62 nsew
rlabel metal3 s 0 11568 800 11688 4 b[5]
port 63 nsew
rlabel metal3 s 1050 12308 1050 12308 4 b[6]
rlabel metal2 s 12282 1588 12282 1588 4 b[7]
rlabel metal3 s 0 16328 800 16448 4 b[8]
port 66 nsew
rlabel metal3 s 1050 15028 1050 15028 4 b[9]
rlabel metal2 s 23690 24021 23690 24021 4 binv
rlabel metal2 s 10994 1588 10994 1588 4 cin
rlabel metal2 s 13570 1520 13570 1520 4 cout
rlabel metal1 s 5290 2312 5290 2312 4 net1
rlabel metal1 s 18412 23698 18412 23698 4 net10
rlabel metal1 s 5014 9928 5014 9928 4 net100
rlabel metal1 s 9292 7174 9292 7174 4 net101
rlabel metal1 s 11178 24786 11178 24786 4 net102
rlabel metal1 s 2185 18734 2185 18734 4 net103
rlabel metal1 s 17296 10166 17296 10166 4 net104
rlabel metal1 s 17526 20434 17526 20434 4 net105
rlabel metal1 s 19504 20978 19504 20978 4 net106
rlabel metal2 s 10994 6596 10994 6596 4 net107
rlabel metal2 s 20010 18564 20010 18564 4 net108
rlabel metal1 s 20792 16218 20792 16218 4 net109
rlabel metal2 s 23120 20910 23120 20910 4 net11
rlabel metal1 s 18722 16218 18722 16218 4 net110
rlabel metal1 s 15594 15470 15594 15470 4 net111
rlabel metal2 s 16238 9180 16238 9180 4 net112
rlabel metal1 s 18630 10778 18630 10778 4 net113
rlabel metal1 s 20286 10098 20286 10098 4 net114
rlabel metal2 s 20930 8092 20930 8092 4 net115
rlabel metal1 s 19366 8466 19366 8466 4 net116
rlabel metal1 s 17802 6766 17802 6766 4 net117
rlabel metal2 s 8694 6052 8694 6052 4 net118
rlabel metal1 s 16054 6290 16054 6290 4 net119
rlabel metal2 s 11914 2992 11914 2992 4 net12
rlabel metal2 s 5566 5508 5566 5508 4 net120
rlabel metal2 s 7314 7684 7314 7684 4 net121
rlabel metal1 s 5566 10030 5566 10030 4 net122
rlabel metal1 s 8142 10030 8142 10030 4 net123
rlabel metal1 s 10488 11866 10488 11866 4 net124
rlabel metal1 s 10120 16218 10120 16218 4 net125
rlabel metal1 s 8326 17646 8326 17646 4 net126
rlabel metal1 s 13616 9010 13616 9010 4 net127
rlabel metal1 s 5290 16660 5290 16660 4 net128
rlabel metal1 s 4922 18394 4922 18394 4 net129
rlabel metal2 s 23580 18258 23580 18258 4 net13
rlabel metal2 s 7130 19652 7130 19652 4 net130
rlabel metal1 s 9430 20434 9430 20434 4 net131
rlabel metal2 s 10626 20060 10626 20060 4 net132
rlabel metal1 s 11960 18258 11960 18258 4 net133
rlabel metal1 s 18170 18394 18170 18394 4 net134
rlabel metal1 s 15318 20434 15318 20434 4 net135
rlabel metal2 s 23518 14382 23518 14382 4 net14
rlabel metal2 s 23690 14960 23690 14960 4 net15
rlabel metal1 s 14794 12818 14794 12818 4 net16
rlabel metal1 s 17802 11798 17802 11798 4 net17
rlabel metal1 s 23506 12716 23506 12716 4 net18
rlabel metal1 s 23414 5882 23414 5882 4 net19
rlabel metal1 s 4508 14246 4508 14246 4 net2
rlabel metal2 s 23518 7854 23518 7854 4 net20
rlabel metal2 s 23506 3876 23506 3876 4 net21
rlabel metal1 s 20470 2618 20470 2618 4 net22
rlabel metal1 s 7406 3094 7406 3094 4 net23
rlabel metal1 s 17434 2618 17434 2618 4 net24
rlabel metal1 s 16008 2550 16008 2550 4 net25
rlabel metal1 s 4692 3094 4692 3094 4 net26
rlabel metal1 s 3697 7378 3697 7378 4 net27
rlabel metal2 s 4968 12206 4968 12206 4 net28
rlabel metal2 s 1610 13022 1610 13022 4 net29
rlabel metal1 s 2185 20774 2185 20774 4 net3
rlabel metal1 s 13294 2618 13294 2618 4 net30
rlabel metal1 s 2185 16966 2185 16966 4 net31
rlabel metal2 s 7406 15538 7406 15538 4 net32
rlabel metal1 s 4830 2958 4830 2958 4 net33
rlabel metal1 s 10810 2618 10810 2618 4 net34
rlabel metal1 s 2185 14246 2185 14246 4 net35
rlabel metal1 s 2185 21658 2185 21658 4 net36
rlabel metal1 s 6808 22610 6808 22610 4 net37
rlabel metal1 s 7958 23766 7958 23766 4 net38
rlabel metal1 s 12006 22746 12006 22746 4 net39
rlabel metal1 s 6440 23086 6440 23086 4 net4
rlabel metal1 s 13368 17170 13368 17170 4 net40
rlabel metal2 s 23598 17595 23598 17595 4 net41
rlabel metal1 s 14812 23834 14812 23834 4 net42
rlabel metal2 s 17618 24208 17618 24208 4 net43
rlabel metal1 s 20700 22746 20700 22746 4 net44
rlabel metal1 s 6256 2550 6256 2550 4 net45
rlabel metal2 s 23518 18734 23518 18734 4 net46
rlabel metal2 s 23580 14994 23580 14994 4 net47
rlabel metal1 s 23506 13804 23506 13804 4 net48
rlabel metal2 s 23230 13566 23230 13566 4 net49
rlabel metal2 s 9338 24208 9338 24208 4 net5
rlabel metal1 s 15479 11118 15479 11118 4 net50
rlabel metal1 s 23506 13362 23506 13362 4 net51
rlabel metal1 s 23672 10642 23672 10642 4 net52
rlabel metal2 s 22954 7990 22954 7990 4 net53
rlabel metal1 s 20636 4590 20636 4590 4 net54
rlabel metal1 s 18704 3026 18704 3026 4 net55
rlabel metal2 s 7360 2550 7360 2550 4 net56
rlabel metal2 s 15042 2924 15042 2924 4 net57
rlabel metal1 s 13046 5678 13046 5678 4 net58
rlabel metal2 s 4554 2822 4554 2822 4 net59
rlabel metal1 s 12512 21998 12512 21998 4 net6
rlabel metal2 s 2622 7582 2622 7582 4 net60
rlabel metal2 s 4830 11968 4830 11968 4 net61
rlabel metal1 s 2185 12682 2185 12682 4 net62
rlabel metal1 s 12604 2618 12604 2618 4 net63
rlabel metal1 s 12581 14314 12581 14314 4 net64
rlabel metal2 s 7038 14994 7038 14994 4 net65
rlabel metal2 s 23046 21522 23046 21522 4 net66
rlabel metal1 s 11500 8466 11500 8466 4 net67
rlabel metal1 s 5290 5134 5290 5134 4 net68
rlabel metal1 s 4922 9486 4922 9486 4 net69
rlabel metal1 s 13018 24582 13018 24582 4 net7
rlabel metal1 s 13478 5542 13478 5542 4 net70
rlabel metal1 s 15916 2414 15916 2414 4 net71
rlabel metal1 s 6900 9010 6900 9010 4 net72
rlabel metal1 s 2185 18258 2185 18258 4 net73
rlabel metal1 s 8786 18394 8786 18394 4 net74
rlabel metal1 s 2185 19346 2185 19346 4 net75
rlabel metal1 s 9246 24786 9246 24786 4 net76
rlabel metal1 s 10350 24786 10350 24786 4 net77
rlabel metal1 s 9936 24786 9936 24786 4 net78
rlabel metal1 s 23184 17646 23184 17646 4 net79
rlabel metal2 s 23874 20230 23874 20230 4 net8
rlabel metal1 s 14398 20026 14398 20026 4 net80
rlabel metal1 s 16238 20026 16238 20026 4 net81
rlabel metal2 s 18814 19652 18814 19652 4 net82
rlabel metal1 s 9890 6630 9890 6630 4 net83
rlabel metal2 s 23230 19142 23230 19142 4 net84
rlabel metal1 s 22793 17170 22793 17170 4 net85
rlabel metal1 s 23644 21522 23644 21522 4 net86
rlabel metal1 s 15042 16218 15042 16218 4 net87
rlabel metal1 s 18170 2414 18170 2414 4 net88
rlabel metal1 s 23552 6766 23552 6766 4 net89
rlabel metal2 s 16882 24378 16882 24378 4 net9
rlabel metal1 s 22793 9554 22793 9554 4 net90
rlabel metal1 s 20884 2414 20884 2414 4 net91
rlabel metal1 s 22793 8942 22793 8942 4 net92
rlabel metal1 s 16606 7174 16606 7174 4 net93
rlabel metal2 s 8602 5865 8602 5865 4 net94
rlabel metal1 s 15962 7242 15962 7242 4 net95
rlabel metal1 s 23506 8500 23506 8500 4 net96
rlabel metal1 s 7314 6630 7314 6630 4 net97
rlabel metal2 s 8050 4794 8050 4794 4 net98
rlabel metal1 s 5152 9350 5152 9350 4 net99
rlabel metal2 s 15502 959 15502 959 4 overflow
rlabel metal3 s 0 8848 800 8968 4 result[0]
port 73 nsew
rlabel metal3 s 1050 17748 1050 17748 4 result[10]
rlabel metal1 s 8464 24650 8464 24650 4 result[11]
rlabel metal3 s 1050 19108 1050 19108 4 result[12]
rlabel metal1 s 9108 24650 9108 24650 4 result[13]
rlabel metal1 s 10534 24650 10534 24650 4 result[14]
rlabel metal1 s 9752 24650 9752 24650 4 result[15]
rlabel metal3 s 23690 17765 23690 17765 4 result[16]
rlabel metal1 s 14260 24650 14260 24650 4 result[17]
rlabel metal1 s 16284 24650 16284 24650 4 result[18]
rlabel metal2 s 23690 19737 23690 19737 4 result[19]
rlabel metal2 s 9706 1520 9706 1520 4 result[1]
rlabel metal2 s 23414 19295 23414 19295 4 result[20]
rlabel metal3 s 23690 17051 23690 17051 4 result[21]
rlabel metal2 s 23690 21233 23690 21233 4 result[22]
rlabel metal1 s 15548 24650 15548 24650 4 result[23]
rlabel metal2 s 18078 1520 18078 1520 4 result[24]
rlabel metal2 s 23690 6749 23690 6749 4 result[25]
rlabel metal2 s 23690 9503 23690 9503 4 result[26]
rlabel metal2 s 20654 1520 20654 1520 4 result[27]
rlabel metal2 s 23690 8857 23690 8857 4 result[28]
rlabel metal2 s 16790 1520 16790 1520 4 result[29]
rlabel metal2 s 8418 1520 8418 1520 4 result[2]
rlabel metal2 s 16146 959 16146 959 4 result[30]
rlabel metal1 s 23552 8330 23552 8330 4 result[31]
rlabel metal2 s 6486 1520 6486 1520 4 result[3]
rlabel metal2 s 7774 1520 7774 1520 4 result[4]
rlabel metal3 s 0 10208 800 10328 4 result[5]
port 100 nsew
rlabel metal3 s 1050 9588 1050 9588 4 result[6]
rlabel metal2 s 9062 1520 9062 1520 4 result[7]
rlabel metal1 s 11040 24650 11040 24650 4 result[8]
rlabel metal3 s 0 18368 800 18488 4 result[9]
port 104 nsew
rlabel metal2 s 23690 4369 23690 4369 4 select[0]
rlabel metal3 s 0 19728 800 19848 4 select[1]
port 106 nsew
rlabel metal2 s 20010 1520 20010 1520 4 zero
flabel metal5 s 1056 22668 24060 22988 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 16956 24060 17276 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 11244 24060 11564 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 5532 24060 5852 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 21648 2128 21968 25072 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 15921 2128 16241 25072 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 10194 2128 10514 25072 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4467 2128 4787 25072 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 22008 24060 22328 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 16296 24060 16616 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 10584 24060 10904 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4872 24060 5192 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 20988 2128 21308 25072 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 15261 2128 15581 25072 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 9534 2128 9854 25072 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3807 2128 4127 25072 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 a[0]
port 3 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 a[10]
port 4 nsew
flabel metal3 s 0 20408 800 20528 0 FreeSans 600 0 0 0 a[11]
port 5 nsew
flabel metal2 s 5814 26516 5870 27316 0 FreeSans 280 90 0 0 a[12]
port 6 nsew
flabel metal2 s 7746 26516 7802 27316 0 FreeSans 280 90 0 0 a[13]
port 7 nsew
flabel metal2 s 12254 26516 12310 27316 0 FreeSans 280 90 0 0 a[14]
port 8 nsew
flabel metal2 s 12898 26516 12954 27316 0 FreeSans 280 90 0 0 a[15]
port 9 nsew
flabel metal3 s 24372 23128 25172 23248 0 FreeSans 600 0 0 0 a[16]
port 10 nsew
flabel metal2 s 16762 26516 16818 27316 0 FreeSans 280 90 0 0 a[17]
port 11 nsew
flabel metal2 s 18050 26516 18106 27316 0 FreeSans 280 90 0 0 a[18]
port 12 nsew
flabel metal3 s 24372 22448 25172 22568 0 FreeSans 600 0 0 0 a[19]
port 13 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 a[1]
port 14 nsew
flabel metal3 s 24372 21768 25172 21888 0 FreeSans 600 0 0 0 a[20]
port 15 nsew
flabel metal3 s 24372 16328 25172 16448 0 FreeSans 600 0 0 0 a[21]
port 16 nsew
flabel metal3 s 24372 14968 25172 15088 0 FreeSans 600 0 0 0 a[22]
port 17 nsew
flabel metal3 s 24372 4768 25172 4888 0 FreeSans 600 0 0 0 a[23]
port 18 nsew
flabel metal3 s 24372 11568 25172 11688 0 FreeSans 600 0 0 0 a[24]
port 19 nsew
flabel metal3 s 24372 12248 25172 12368 0 FreeSans 600 0 0 0 a[25]
port 20 nsew
flabel metal3 s 24372 5448 25172 5568 0 FreeSans 600 0 0 0 a[26]
port 21 nsew
flabel metal3 s 24372 6128 25172 6248 0 FreeSans 600 0 0 0 a[27]
port 22 nsew
flabel metal3 s 24372 2728 25172 2848 0 FreeSans 600 0 0 0 a[28]
port 23 nsew
flabel metal2 s 21270 0 21326 800 0 FreeSans 280 90 0 0 a[29]
port 24 nsew
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 a[2]
port 25 nsew
flabel metal2 s 18694 0 18750 800 0 FreeSans 280 90 0 0 a[30]
port 26 nsew
flabel metal2 s 14830 0 14886 800 0 FreeSans 280 90 0 0 a[31]
port 27 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 a[3]
port 28 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 a[4]
port 29 nsew
flabel metal3 s 0 10888 800 11008 0 FreeSans 600 0 0 0 a[5]
port 30 nsew
flabel metal3 s 400 12988 400 12988 0 FreeSans 600 0 0 0 a[6]
flabel metal2 s 12898 0 12954 800 0 FreeSans 280 90 0 0 a[7]
port 32 nsew
flabel metal3 s 400 17068 400 17068 0 FreeSans 600 0 0 0 a[8]
flabel metal3 s 400 15708 400 15708 0 FreeSans 600 0 0 0 a[9]
flabel metal3 s 24372 24488 25172 24608 0 FreeSans 600 0 0 0 ainv
port 35 nsew
flabel metal2 s 10322 0 10378 800 0 FreeSans 280 90 0 0 b[0]
port 36 nsew
flabel metal3 s 400 14348 400 14348 0 FreeSans 600 0 0 0 b[10]
flabel metal3 s 400 21148 400 21148 0 FreeSans 600 0 0 0 b[11]
flabel metal2 s 6458 26516 6514 27316 0 FreeSans 280 90 0 0 b[12]
port 39 nsew
flabel metal2 s 7102 26516 7158 27316 0 FreeSans 280 90 0 0 b[13]
port 40 nsew
flabel metal2 s 11610 26516 11666 27316 0 FreeSans 280 90 0 0 b[14]
port 41 nsew
flabel metal2 s 13542 26516 13598 27316 0 FreeSans 280 90 0 0 b[15]
port 42 nsew
flabel metal3 s 24372 18368 25172 18488 0 FreeSans 600 0 0 0 b[16]
port 43 nsew
flabel metal2 s 14830 26516 14886 27316 0 FreeSans 280 90 0 0 b[17]
port 44 nsew
flabel metal2 s 17406 26516 17462 27316 0 FreeSans 280 90 0 0 b[18]
port 45 nsew
flabel metal2 s 20626 26516 20682 27316 0 FreeSans 280 90 0 0 b[19]
port 46 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 b[1]
port 47 nsew
flabel metal3 s 24372 20408 25172 20528 0 FreeSans 600 0 0 0 b[20]
port 48 nsew
flabel metal3 s 24372 15648 25172 15768 0 FreeSans 600 0 0 0 b[21]
port 49 nsew
flabel metal3 s 24372 14288 25172 14408 0 FreeSans 600 0 0 0 b[22]
port 50 nsew
flabel metal3 s 24372 13608 25172 13728 0 FreeSans 600 0 0 0 b[23]
port 51 nsew
flabel metal3 s 24372 10888 25172 11008 0 FreeSans 600 0 0 0 b[24]
port 52 nsew
flabel metal3 s 24372 12928 25172 13048 0 FreeSans 600 0 0 0 b[25]
port 53 nsew
flabel metal3 s 24372 10208 25172 10328 0 FreeSans 600 0 0 0 b[26]
port 54 nsew
flabel metal3 s 24372 7488 25172 7608 0 FreeSans 600 0 0 0 b[27]
port 55 nsew
flabel metal3 s 24372 3408 25172 3528 0 FreeSans 600 0 0 0 b[28]
port 56 nsew
flabel metal2 s 19338 0 19394 800 0 FreeSans 280 90 0 0 b[29]
port 57 nsew
flabel metal2 s 7102 0 7158 800 0 FreeSans 280 90 0 0 b[2]
port 58 nsew
flabel metal2 s 17406 0 17462 800 0 FreeSans 280 90 0 0 b[30]
port 59 nsew
flabel metal2 s 14186 0 14242 800 0 FreeSans 280 90 0 0 b[31]
port 60 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 b[3]
port 61 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 b[4]
flabel metal3 s 400 11628 400 11628 0 FreeSans 600 0 0 0 b[5]
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 b[6]
port 64 nsew
flabel metal2 s 12254 0 12310 800 0 FreeSans 280 90 0 0 b[7]
port 65 nsew
flabel metal3 s 400 16388 400 16388 0 FreeSans 600 0 0 0 b[8]
flabel metal3 s 0 14968 800 15088 0 FreeSans 600 0 0 0 b[9]
port 67 nsew
flabel metal3 s 24372 23808 25172 23928 0 FreeSans 600 0 0 0 binv
port 68 nsew
flabel metal2 s 10966 0 11022 800 0 FreeSans 280 90 0 0 cin
port 69 nsew
flabel metal2 s 13542 0 13598 800 0 FreeSans 280 90 0 0 cout
port 70 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 fake_clk
port 71 nsew
flabel metal2 s 15474 0 15530 800 0 FreeSans 280 90 0 0 overflow
port 72 nsew
flabel metal3 s 400 8908 400 8908 0 FreeSans 600 0 0 0 result[0]
flabel metal3 s 0 17688 800 17808 0 FreeSans 600 0 0 0 result[10]
port 74 nsew
flabel metal2 s 8390 26516 8446 27316 0 FreeSans 280 90 0 0 result[11]
port 75 nsew
flabel metal3 s 0 19048 800 19168 0 FreeSans 600 0 0 0 result[12]
port 76 nsew
flabel metal2 s 9034 26516 9090 27316 0 FreeSans 280 90 0 0 result[13]
port 77 nsew
flabel metal2 s 10322 26516 10378 27316 0 FreeSans 280 90 0 0 result[14]
port 78 nsew
flabel metal2 s 9678 26516 9734 27316 0 FreeSans 280 90 0 0 result[15]
port 79 nsew
flabel metal3 s 24372 17688 25172 17808 0 FreeSans 600 0 0 0 result[16]
port 80 nsew
flabel metal2 s 14186 26516 14242 27316 0 FreeSans 280 90 0 0 result[17]
port 81 nsew
flabel metal2 s 16118 26516 16174 27316 0 FreeSans 280 90 0 0 result[18]
port 82 nsew
flabel metal3 s 24372 19728 25172 19848 0 FreeSans 600 0 0 0 result[19]
port 83 nsew
flabel metal2 s 9678 0 9734 800 0 FreeSans 280 90 0 0 result[1]
port 84 nsew
flabel metal3 s 24372 19048 25172 19168 0 FreeSans 600 0 0 0 result[20]
port 85 nsew
flabel metal3 s 24372 17008 25172 17128 0 FreeSans 600 0 0 0 result[21]
port 86 nsew
flabel metal3 s 24372 21088 25172 21208 0 FreeSans 600 0 0 0 result[22]
port 87 nsew
flabel metal2 s 15474 26516 15530 27316 0 FreeSans 280 90 0 0 result[23]
port 88 nsew
flabel metal2 s 18050 0 18106 800 0 FreeSans 280 90 0 0 result[24]
port 89 nsew
flabel metal3 s 24372 6808 25172 6928 0 FreeSans 600 0 0 0 result[25]
port 90 nsew
flabel metal3 s 24372 9528 25172 9648 0 FreeSans 600 0 0 0 result[26]
port 91 nsew
flabel metal2 s 20626 0 20682 800 0 FreeSans 280 90 0 0 result[27]
port 92 nsew
flabel metal3 s 24372 8848 25172 8968 0 FreeSans 600 0 0 0 result[28]
port 93 nsew
flabel metal2 s 16762 0 16818 800 0 FreeSans 280 90 0 0 result[29]
port 94 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 result[2]
port 95 nsew
flabel metal2 s 16118 0 16174 800 0 FreeSans 280 90 0 0 result[30]
port 96 nsew
flabel metal3 s 24372 8168 25172 8288 0 FreeSans 600 0 0 0 result[31]
port 97 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 result[3]
port 98 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 result[4]
port 99 nsew
flabel metal3 s 400 10268 400 10268 0 FreeSans 600 0 0 0 result[5]
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 result[6]
port 101 nsew
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 result[7]
port 102 nsew
flabel metal2 s 10966 26516 11022 27316 0 FreeSans 280 90 0 0 result[8]
port 103 nsew
flabel metal3 s 400 18428 400 18428 0 FreeSans 600 0 0 0 result[9]
flabel metal3 s 24372 4088 25172 4208 0 FreeSans 600 0 0 0 select[0]
port 105 nsew
flabel metal3 s 400 19788 400 19788 0 FreeSans 600 0 0 0 select[1]
flabel metal2 s 19982 0 20038 800 0 FreeSans 280 90 0 0 zero
port 107 nsew
<< properties >>
string FIXED_BBOX 0 0 25172 27316
<< end >>
