VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO n_bit_alu
  CLASS BLOCK ;
  FOREIGN n_bit_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 117.340 BY 128.060 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.300 10.640 22.900 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.865 10.640 49.465 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.430 10.640 76.030 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.995 10.640 102.595 117.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.640 112.020 28.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 53.160 112.020 54.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 79.680 112.020 81.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 106.200 112.020 107.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.000 10.640 19.600 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.565 10.640 46.165 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.130 10.640 72.730 117.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.695 10.640 99.295 117.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 23.340 112.020 24.940 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 49.860 112.020 51.460 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.380 112.020 77.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 102.900 112.020 104.500 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 124.060 26.130 128.060 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 124.060 42.230 128.060 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 124.060 45.450 128.060 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 124.060 55.110 128.060 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 124.060 77.650 128.060 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 124.060 67.990 128.060 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 124.060 93.750 128.060 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 102.040 117.340 102.640 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 98.640 117.340 99.240 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 78.240 117.340 78.840 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 95.240 117.340 95.840 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 61.240 117.340 61.840 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 57.840 117.340 58.440 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 71.440 117.340 72.040 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 23.840 117.340 24.440 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 27.240 117.340 27.840 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 20.440 117.340 21.040 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END a[9]
  PIN ainv
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END ainv
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 124.060 22.910 128.060 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 124.060 32.570 128.060 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 124.060 48.670 128.060 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 124.060 51.890 128.060 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 124.060 74.430 128.060 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 124.060 64.770 128.060 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 124.060 87.310 128.060 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 124.060 96.970 128.060 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 91.840 117.340 92.440 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 74.840 117.340 75.440 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 81.640 117.340 82.240 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 68.040 117.340 68.640 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 54.440 117.340 55.040 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 64.640 117.340 65.240 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 51.040 117.340 51.640 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 34.040 117.340 34.640 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END b[9]
  PIN binv
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END binv
  PIN cin
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END cin
  PIN cout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END cout
  PIN fake_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END fake_clk
  PIN overflow
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END overflow
  PIN result[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END result[0]
  PIN result[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END result[10]
  PIN result[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END result[11]
  PIN result[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END result[12]
  PIN result[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 124.060 35.790 128.060 ;
    END
  END result[13]
  PIN result[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.730 124.060 39.010 128.060 ;
    END
  END result[14]
  PIN result[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END result[15]
  PIN result[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 124.060 90.530 128.060 ;
    END
  END result[16]
  PIN result[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.270 124.060 61.550 128.060 ;
    END
  END result[17]
  PIN result[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 124.060 71.210 128.060 ;
    END
  END result[18]
  PIN result[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 124.060 80.870 128.060 ;
    END
  END result[19]
  PIN result[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END result[1]
  PIN result[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 124.060 84.090 128.060 ;
    END
  END result[20]
  PIN result[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 88.440 117.340 89.040 ;
    END
  END result[21]
  PIN result[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 85.040 117.340 85.640 ;
    END
  END result[22]
  PIN result[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.050 124.060 58.330 128.060 ;
    END
  END result[23]
  PIN result[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END result[24]
  PIN result[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 30.640 117.340 31.240 ;
    END
  END result[25]
  PIN result[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 47.640 117.340 48.240 ;
    END
  END result[26]
  PIN result[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 37.440 117.340 38.040 ;
    END
  END result[27]
  PIN result[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 40.840 117.340 41.440 ;
    END
  END result[28]
  PIN result[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END result[29]
  PIN result[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END result[2]
  PIN result[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END result[30]
  PIN result[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 113.340 44.240 117.340 44.840 ;
    END
  END result[31]
  PIN result[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END result[7]
  PIN result[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END result[8]
  PIN result[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END result[9]
  PIN select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END select[0]
  PIN select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END select[1]
  PIN zero
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END zero
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 111.970 117.150 ;
      LAYER li1 ;
        RECT 5.520 10.795 111.780 117.045 ;
      LAYER met1 ;
        RECT 4.210 10.640 111.780 117.200 ;
      LAYER met2 ;
        RECT 4.230 123.780 22.350 124.850 ;
        RECT 23.190 123.780 25.570 124.850 ;
        RECT 26.410 123.780 32.010 124.850 ;
        RECT 32.850 123.780 35.230 124.850 ;
        RECT 36.070 123.780 38.450 124.850 ;
        RECT 39.290 123.780 41.670 124.850 ;
        RECT 42.510 123.780 44.890 124.850 ;
        RECT 45.730 123.780 48.110 124.850 ;
        RECT 48.950 123.780 51.330 124.850 ;
        RECT 52.170 123.780 54.550 124.850 ;
        RECT 55.390 123.780 57.770 124.850 ;
        RECT 58.610 123.780 60.990 124.850 ;
        RECT 61.830 123.780 64.210 124.850 ;
        RECT 65.050 123.780 67.430 124.850 ;
        RECT 68.270 123.780 70.650 124.850 ;
        RECT 71.490 123.780 73.870 124.850 ;
        RECT 74.710 123.780 77.090 124.850 ;
        RECT 77.930 123.780 80.310 124.850 ;
        RECT 81.150 123.780 83.530 124.850 ;
        RECT 84.370 123.780 86.750 124.850 ;
        RECT 87.590 123.780 89.970 124.850 ;
        RECT 90.810 123.780 93.190 124.850 ;
        RECT 94.030 123.780 96.410 124.850 ;
        RECT 97.250 123.780 110.310 124.850 ;
        RECT 4.230 4.280 110.310 123.780 ;
        RECT 4.230 3.670 15.910 4.280 ;
        RECT 16.750 3.670 19.130 4.280 ;
        RECT 19.970 3.670 22.350 4.280 ;
        RECT 23.190 3.670 25.570 4.280 ;
        RECT 26.410 3.670 28.790 4.280 ;
        RECT 29.630 3.670 32.010 4.280 ;
        RECT 32.850 3.670 35.230 4.280 ;
        RECT 36.070 3.670 38.450 4.280 ;
        RECT 39.290 3.670 41.670 4.280 ;
        RECT 42.510 3.670 44.890 4.280 ;
        RECT 45.730 3.670 48.110 4.280 ;
        RECT 48.950 3.670 51.330 4.280 ;
        RECT 52.170 3.670 54.550 4.280 ;
        RECT 55.390 3.670 57.770 4.280 ;
        RECT 58.610 3.670 60.990 4.280 ;
        RECT 61.830 3.670 64.210 4.280 ;
        RECT 65.050 3.670 67.430 4.280 ;
        RECT 68.270 3.670 70.650 4.280 ;
        RECT 71.490 3.670 73.870 4.280 ;
        RECT 74.710 3.670 77.090 4.280 ;
        RECT 77.930 3.670 80.310 4.280 ;
        RECT 81.150 3.670 83.530 4.280 ;
        RECT 84.370 3.670 86.750 4.280 ;
        RECT 87.590 3.670 89.970 4.280 ;
        RECT 90.810 3.670 93.190 4.280 ;
        RECT 94.030 3.670 96.410 4.280 ;
        RECT 97.250 3.670 99.630 4.280 ;
        RECT 100.470 3.670 110.310 4.280 ;
      LAYER met3 ;
        RECT 3.990 113.240 113.340 117.125 ;
        RECT 4.400 111.840 113.340 113.240 ;
        RECT 3.990 109.840 113.340 111.840 ;
        RECT 4.400 108.440 113.340 109.840 ;
        RECT 3.990 106.440 113.340 108.440 ;
        RECT 4.400 105.040 113.340 106.440 ;
        RECT 3.990 103.040 113.340 105.040 ;
        RECT 4.400 101.640 112.940 103.040 ;
        RECT 3.990 99.640 113.340 101.640 ;
        RECT 4.400 98.240 112.940 99.640 ;
        RECT 3.990 96.240 113.340 98.240 ;
        RECT 4.400 94.840 112.940 96.240 ;
        RECT 3.990 92.840 113.340 94.840 ;
        RECT 4.400 91.440 112.940 92.840 ;
        RECT 3.990 89.440 113.340 91.440 ;
        RECT 4.400 88.040 112.940 89.440 ;
        RECT 3.990 86.040 113.340 88.040 ;
        RECT 4.400 84.640 112.940 86.040 ;
        RECT 3.990 82.640 113.340 84.640 ;
        RECT 4.400 81.240 112.940 82.640 ;
        RECT 3.990 79.240 113.340 81.240 ;
        RECT 4.400 77.840 112.940 79.240 ;
        RECT 3.990 75.840 113.340 77.840 ;
        RECT 4.400 74.440 112.940 75.840 ;
        RECT 3.990 72.440 113.340 74.440 ;
        RECT 4.400 71.040 112.940 72.440 ;
        RECT 3.990 69.040 113.340 71.040 ;
        RECT 4.400 67.640 112.940 69.040 ;
        RECT 3.990 65.640 113.340 67.640 ;
        RECT 4.400 64.240 112.940 65.640 ;
        RECT 3.990 62.240 113.340 64.240 ;
        RECT 4.400 60.840 112.940 62.240 ;
        RECT 3.990 58.840 113.340 60.840 ;
        RECT 4.400 57.440 112.940 58.840 ;
        RECT 3.990 55.440 113.340 57.440 ;
        RECT 4.400 54.040 112.940 55.440 ;
        RECT 3.990 52.040 113.340 54.040 ;
        RECT 4.400 50.640 112.940 52.040 ;
        RECT 3.990 48.640 113.340 50.640 ;
        RECT 4.400 47.240 112.940 48.640 ;
        RECT 3.990 45.240 113.340 47.240 ;
        RECT 4.400 43.840 112.940 45.240 ;
        RECT 3.990 41.840 113.340 43.840 ;
        RECT 4.400 40.440 112.940 41.840 ;
        RECT 3.990 38.440 113.340 40.440 ;
        RECT 4.400 37.040 112.940 38.440 ;
        RECT 3.990 35.040 113.340 37.040 ;
        RECT 4.400 33.640 112.940 35.040 ;
        RECT 3.990 31.640 113.340 33.640 ;
        RECT 4.400 30.240 112.940 31.640 ;
        RECT 3.990 28.240 113.340 30.240 ;
        RECT 4.400 26.840 112.940 28.240 ;
        RECT 3.990 24.840 113.340 26.840 ;
        RECT 4.400 23.440 112.940 24.840 ;
        RECT 3.990 21.440 113.340 23.440 ;
        RECT 4.400 20.040 112.940 21.440 ;
        RECT 3.990 18.040 113.340 20.040 ;
        RECT 4.400 16.640 113.340 18.040 ;
        RECT 3.990 10.715 113.340 16.640 ;
  END
END n_bit_alu
END LIBRARY

