module n_bit_alu (ainv,
    binv,
    cin,
    cout,
    fake_clk,
    overflow,
    zero,
    a,
    b,
    result,
    select);
 input ainv;
 input binv;
 input cin;
 output cout;
 input fake_clk;
 output overflow;
 output zero;
 input [31:0] a;
 input [31:0] b;
 output [31:0] result;
 input [1:0] select;

 wire _0030_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0090_;
 wire _0094_;
 wire _0105_;
 wire _0108_;
 wire _0111_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0131_;
 wire _0146_;
 wire _0152_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0172_;
 wire _0176_;
 wire _0178_;
 wire _0187_;
 wire _0193_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0213_;
 wire _0217_;
 wire _0228_;
 wire _0234_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0254_;
 wire _0258_;
 wire _0269_;
 wire _0275_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0295_;
 wire _0299_;
 wire _0310_;
 wire _0316_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0336_;
 wire _0340_;
 wire _0351_;
 wire _0357_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0377_;
 wire _0381_;
 wire _0392_;
 wire _0398_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0418_;
 wire _0422_;
 wire _0433_;
 wire _0439_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0459_;
 wire _0463_;
 wire _0474_;
 wire _0480_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0500_;
 wire _0504_;
 wire _0515_;
 wire _0521_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0541_;
 wire _0545_;
 wire _0556_;
 wire _0562_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0582_;
 wire _0586_;
 wire _0597_;
 wire _0603_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0623_;
 wire _0627_;
 wire _0638_;
 wire _0644_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0664_;
 wire _0668_;
 wire _0679_;
 wire _0685_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0705_;
 wire _0709_;
 wire _0720_;
 wire _0726_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0746_;
 wire _0750_;
 wire _0761_;
 wire _0767_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0787_;
 wire _0791_;
 wire _0802_;
 wire _0808_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0828_;
 wire _0832_;
 wire _0843_;
 wire _0849_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0869_;
 wire _0873_;
 wire _0884_;
 wire _0890_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0910_;
 wire _0914_;
 wire _0925_;
 wire _0931_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0951_;
 wire _0955_;
 wire _0966_;
 wire _0972_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0992_;
 wire _0996_;
 wire _1007_;
 wire _1013_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1033_;
 wire _1037_;
 wire _1048_;
 wire _1054_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1074_;
 wire _1078_;
 wire _1089_;
 wire _1095_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1115_;
 wire _1119_;
 wire _1130_;
 wire _1136_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1156_;
 wire _1160_;
 wire _1171_;
 wire _1177_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1197_;
 wire _1201_;
 wire _1212_;
 wire _1218_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1238_;
 wire _1242_;
 wire _1253_;
 wire _1259_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1279_;
 wire _1283_;
 wire _1294_;
 wire _1300_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1320_;
 wire _1324_;
 wire _1335_;
 wire _1341_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1361_;
 wire _1365_;
 wire _1376_;
 wire _1382_;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net129;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;

 sky130_fd_sc_hd__nor4_1 _1388_ (.A(_0050_),
    .B(_0053_),
    .C(_0056_),
    .D(_0057_),
    .Y(_0032_));
 sky130_fd_sc_hd__nor4_4 _1389_ (.A(_0060_),
    .B(_0061_),
    .C(_0063_),
    .D(_0067_),
    .Y(_0033_));
 sky130_fd_sc_hd__nor4_1 _1390_ (.A(_0054_),
    .B(_0065_),
    .C(_0069_),
    .D(_0072_),
    .Y(_0034_));
 sky130_fd_sc_hd__nor4_1 _1391_ (.A(_0073_),
    .B(_0045_),
    .C(_0047_),
    .D(_0048_),
    .Y(_0035_));
 sky130_fd_sc_hd__nand4_1 _1392_ (.A(_0033_),
    .B(_0032_),
    .C(_0034_),
    .D(net106),
    .Y(_0036_));
 sky130_fd_sc_hd__nor4_1 _1393_ (.A(_0051_),
    .B(_0052_),
    .C(_0055_),
    .D(_0058_),
    .Y(_0037_));
 sky130_fd_sc_hd__nor4_2 _1394_ (.A(_0059_),
    .B(_0062_),
    .C(_0066_),
    .D(_0064_),
    .Y(_0038_));
 sky130_fd_sc_hd__nor4_4 _1395_ (.A(_0071_),
    .B(_0068_),
    .C(_0070_),
    .D(_0043_),
    .Y(_0039_));
 sky130_fd_sc_hd__nor4_1 _1396_ (.A(_0074_),
    .B(_0044_),
    .C(_0046_),
    .D(_0049_),
    .Y(_0040_));
 sky130_fd_sc_hd__nand4_1 _1397_ (.A(_0039_),
    .B(_0038_),
    .C(_0037_),
    .D(net105),
    .Y(_0041_));
 sky130_fd_sc_hd__nor2_1 _1398_ (.A(_0036_),
    .B(_0041_),
    .Y(net104));
 sky130_fd_sc_hd__xor2_1 _1399_ (.A(net70),
    .B(_0030_),
    .X(net71));
 sky130_fd_sc_hd__inv_1 _1400_ (.A(net1),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_1 _1401_ (.A(net34),
    .Y(_0080_));
 sky130_fd_sc_hd__and2_0 _1402_ (.A(_0084_),
    .B(_0082_),
    .X(_0081_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1403_ (.A(_0084_),
    .SLEEP(_0082_),
    .X(_0085_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1404_ (.A(_0086_),
    .SLEEP(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__and2_0 _1405_ (.A(_0084_),
    .B(_0082_),
    .X(_0086_));
 sky130_fd_sc_hd__xor2_2 _1406_ (.A(_0084_),
    .B(_0082_),
    .X(_0090_));
 sky130_fd_sc_hd__and2_0 _1407_ (.A(_0090_),
    .B(net67),
    .X(_0087_));
 sky130_fd_sc_hd__xor2_1 _1408_ (.A(net67),
    .B(_0090_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_4 _1409_ (.A0(net1),
    .A1(_0079_),
    .S(net124),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_4 _1410_ (.A0(net34),
    .A1(_0080_),
    .S(net120),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_4 _1411_ (.A0(_0094_),
    .A1(_0108_),
    .S(net111),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_4 _1412_ (.A0(_0111_),
    .A1(_0105_),
    .S(net107),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1413_ (.A0(_0081_),
    .A1(_0085_),
    .S(net111),
    .X(_0111_));
 sky130_fd_sc_hd__inv_1 _1414_ (.A(net25),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_1 _1415_ (.A(net58),
    .Y(_0121_));
 sky130_fd_sc_hd__and2_0 _1416_ (.A(_0125_),
    .B(_0123_),
    .X(_0122_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1417_ (.A(_0125_),
    .SLEEP(_0123_),
    .X(_0126_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1418_ (.A(_0127_),
    .SLEEP(_0128_),
    .X(net70));
 sky130_fd_sc_hd__and2_0 _1419_ (.A(_0125_),
    .B(_0123_),
    .X(_0127_));
 sky130_fd_sc_hd__xor2_1 _1420_ (.A(_0125_),
    .B(_0123_),
    .X(_0131_));
 sky130_fd_sc_hd__and2_0 _1421_ (.A(_0030_),
    .B(_0131_),
    .X(_0128_));
 sky130_fd_sc_hd__xor2_1 _1422_ (.A(_0030_),
    .B(_0131_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1423_ (.A0(net25),
    .A1(_0120_),
    .S(net160),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1424_ (.A0(net58),
    .A1(_0121_),
    .S(net159),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_4 _1425_ (.A0(_0108_),
    .A1(net150),
    .S(net113),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_4 _1426_ (.A0(_0152_),
    .A1(_0146_),
    .S(net107),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1427_ (.A0(_0122_),
    .A1(_0126_),
    .S(net113),
    .X(_0152_));
 sky130_fd_sc_hd__inv_1 _1428_ (.A(net2),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_1 _1429_ (.A(net35),
    .Y(_0162_));
 sky130_fd_sc_hd__and2_0 _1430_ (.A(_0166_),
    .B(_0164_),
    .X(_0163_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1431_ (.A(_0166_),
    .SLEEP(_0164_),
    .X(_0167_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1432_ (.A(_0168_),
    .SLEEP(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_0 _1433_ (.A(_0166_),
    .B(_0164_),
    .X(_0168_));
 sky130_fd_sc_hd__xor2_1 _1434_ (.A(_0166_),
    .B(_0164_),
    .X(_0172_));
 sky130_fd_sc_hd__and2_4 _1435_ (.A(_0178_),
    .B(_0172_),
    .X(_0169_));
 sky130_fd_sc_hd__xor2_1 _1436_ (.A(_0178_),
    .B(_0172_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _1437_ (.A0(net2),
    .A1(_0161_),
    .S(net126),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(net35),
    .A1(_0162_),
    .S(net122),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(_0176_),
    .A1(net151),
    .S(net115),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(_0193_),
    .A1(_0187_),
    .S(net109),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(_0163_),
    .A1(_0167_),
    .S(net115),
    .X(_0193_));
 sky130_fd_sc_hd__inv_1 _1442_ (.A(net3),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_1 _1443_ (.A(net36),
    .Y(_0203_));
 sky130_fd_sc_hd__and2_0 _1444_ (.A(_0207_),
    .B(_0205_),
    .X(_0204_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1445_ (.A(_0207_),
    .SLEEP(_0205_),
    .X(_0208_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1446_ (.A(_0209_),
    .SLEEP(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__and2_0 _1447_ (.A(_0207_),
    .B(_0205_),
    .X(_0209_));
 sky130_fd_sc_hd__xor2_1 _1448_ (.A(_0207_),
    .B(_0205_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_4 _1449_ (.A(_0170_),
    .B(_0213_),
    .X(_0210_));
 sky130_fd_sc_hd__xor2_1 _1450_ (.A(_0170_),
    .B(_0213_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(net3),
    .A1(_0202_),
    .S(net126),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(net36),
    .A1(_0203_),
    .S(net122),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _1453_ (.A0(_0217_),
    .A1(net152),
    .S(net115),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _1454_ (.A0(_0234_),
    .A1(_0228_),
    .S(net109),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _1455_ (.A0(_0204_),
    .A1(_0208_),
    .S(net115),
    .X(_0234_));
 sky130_fd_sc_hd__inv_1 _1456_ (.A(net4),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_1 _1457_ (.A(net37),
    .Y(_0244_));
 sky130_fd_sc_hd__and2_0 _1458_ (.A(_0248_),
    .B(_0246_),
    .X(_0245_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1459_ (.A(_0248_),
    .SLEEP(_0246_),
    .X(_0249_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1460_ (.A(_0250_),
    .SLEEP(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__and2_0 _1461_ (.A(_0248_),
    .B(_0246_),
    .X(_0250_));
 sky130_fd_sc_hd__xor2_1 _1462_ (.A(_0248_),
    .B(_0246_),
    .X(_0254_));
 sky130_fd_sc_hd__and2_4 _1463_ (.A(_0211_),
    .B(_0254_),
    .X(_0251_));
 sky130_fd_sc_hd__xor2_1 _1464_ (.A(_0211_),
    .B(_0254_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(net4),
    .A1(_0243_),
    .S(net126),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _1466_ (.A0(net37),
    .A1(_0244_),
    .S(net122),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(_0258_),
    .A1(net153),
    .S(net116),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(_0275_),
    .A1(_0269_),
    .S(net109),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _1469_ (.A0(_0245_),
    .A1(_0249_),
    .S(net116),
    .X(_0275_));
 sky130_fd_sc_hd__inv_1 _1470_ (.A(net5),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_1 _1471_ (.A(net38),
    .Y(_0285_));
 sky130_fd_sc_hd__and2_0 _1472_ (.A(_0289_),
    .B(_0287_),
    .X(_0286_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1473_ (.A(_0289_),
    .SLEEP(_0287_),
    .X(_0290_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1474_ (.A(_0291_),
    .SLEEP(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__and2_0 _1475_ (.A(_0289_),
    .B(_0287_),
    .X(_0291_));
 sky130_fd_sc_hd__xor2_1 _1476_ (.A(_0289_),
    .B(_0287_),
    .X(_0295_));
 sky130_fd_sc_hd__and2_0 _1477_ (.A(_0295_),
    .B(_0252_),
    .X(_0292_));
 sky130_fd_sc_hd__xor2_1 _1478_ (.A(_0252_),
    .B(_0295_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _1479_ (.A0(net5),
    .A1(_0284_),
    .S(net126),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _1480_ (.A0(net38),
    .A1(_0285_),
    .S(net122),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _1481_ (.A0(_0299_),
    .A1(net154),
    .S(net116),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _1482_ (.A0(_0316_),
    .A1(_0310_),
    .S(net109),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(_0286_),
    .A1(_0290_),
    .S(net116),
    .X(_0316_));
 sky130_fd_sc_hd__inv_1 _1484_ (.A(net6),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_1 _1485_ (.A(net39),
    .Y(_0326_));
 sky130_fd_sc_hd__and2_0 _1486_ (.A(_0330_),
    .B(_0328_),
    .X(_0327_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1487_ (.A(_0330_),
    .SLEEP(_0328_),
    .X(_0331_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1488_ (.A(_0332_),
    .SLEEP(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__and2_0 _1489_ (.A(_0330_),
    .B(_0328_),
    .X(_0332_));
 sky130_fd_sc_hd__xor2_1 _1490_ (.A(_0330_),
    .B(_0328_),
    .X(_0336_));
 sky130_fd_sc_hd__and2_4 _1491_ (.A(_0293_),
    .B(_0336_),
    .X(_0333_));
 sky130_fd_sc_hd__xor2_1 _1492_ (.A(_0293_),
    .B(_0336_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(net6),
    .A1(_0325_),
    .S(net126),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _1494_ (.A0(net39),
    .A1(_0326_),
    .S(net122),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(_0340_),
    .A1(net155),
    .S(net116),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _1496_ (.A0(_0357_),
    .A1(_0351_),
    .S(net109),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(_0327_),
    .A1(_0331_),
    .S(net116),
    .X(_0357_));
 sky130_fd_sc_hd__inv_1 _1498_ (.A(net7),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_1 _1499_ (.A(net40),
    .Y(_0367_));
 sky130_fd_sc_hd__and2_0 _1500_ (.A(_0371_),
    .B(_0369_),
    .X(_0368_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1501_ (.A(_0371_),
    .SLEEP(_0369_),
    .X(_0372_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1502_ (.A(_0373_),
    .SLEEP(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__and2_0 _1503_ (.A(_0371_),
    .B(_0369_),
    .X(_0373_));
 sky130_fd_sc_hd__xor2_1 _1504_ (.A(_0371_),
    .B(_0369_),
    .X(_0377_));
 sky130_fd_sc_hd__and2_4 _1505_ (.A(_0334_),
    .B(_0377_),
    .X(_0374_));
 sky130_fd_sc_hd__xor2_1 _1506_ (.A(_0334_),
    .B(_0377_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(net7),
    .A1(_0366_),
    .S(net126),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _1508_ (.A0(net40),
    .A1(_0367_),
    .S(net122),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _1509_ (.A0(_0381_),
    .A1(net156),
    .S(net115),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(_0398_),
    .A1(_0392_),
    .S(net109),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1511_ (.A0(_0368_),
    .A1(_0372_),
    .S(net115),
    .X(_0398_));
 sky130_fd_sc_hd__inv_1 _1512_ (.A(net8),
    .Y(_0407_));
 sky130_fd_sc_hd__inv_1 _1513_ (.A(net41),
    .Y(_0408_));
 sky130_fd_sc_hd__and2_0 _1514_ (.A(_0412_),
    .B(_0410_),
    .X(_0409_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1515_ (.A(_0412_),
    .SLEEP(_0410_),
    .X(_0413_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1516_ (.A(_0414_),
    .SLEEP(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__and2_0 _1517_ (.A(_0412_),
    .B(_0410_),
    .X(_0414_));
 sky130_fd_sc_hd__xor2_1 _1518_ (.A(_0412_),
    .B(_0410_),
    .X(_0418_));
 sky130_fd_sc_hd__and2_4 _1519_ (.A(_0375_),
    .B(_0418_),
    .X(_0415_));
 sky130_fd_sc_hd__xor2_1 _1520_ (.A(_0375_),
    .B(_0418_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _1521_ (.A0(net8),
    .A1(_0407_),
    .S(net126),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _1522_ (.A0(net41),
    .A1(_0408_),
    .S(net122),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _1523_ (.A0(_0422_),
    .A1(net157),
    .S(net117),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _1524_ (.A0(_0439_),
    .A1(_0433_),
    .S(net109),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(_0409_),
    .A1(_0413_),
    .S(net117),
    .X(_0439_));
 sky130_fd_sc_hd__inv_1 _1526_ (.A(net9),
    .Y(_0448_));
 sky130_fd_sc_hd__inv_1 _1527_ (.A(net42),
    .Y(_0449_));
 sky130_fd_sc_hd__and2_0 _1528_ (.A(_0453_),
    .B(_0451_),
    .X(_0450_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1529_ (.A(_0453_),
    .SLEEP(_0451_),
    .X(_0454_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1530_ (.A(_0455_),
    .SLEEP(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__and2_0 _1531_ (.A(_0453_),
    .B(_0451_),
    .X(_0455_));
 sky130_fd_sc_hd__xor2_1 _1532_ (.A(_0453_),
    .B(_0451_),
    .X(_0459_));
 sky130_fd_sc_hd__and2_4 _1533_ (.A(_0416_),
    .B(_0459_),
    .X(_0456_));
 sky130_fd_sc_hd__xor2_1 _1534_ (.A(_0416_),
    .B(_0459_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _1535_ (.A0(net9),
    .A1(_0448_),
    .S(net126),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(net42),
    .A1(_0449_),
    .S(net122),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _1537_ (.A0(_0463_),
    .A1(net158),
    .S(net117),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1538_ (.A0(_0480_),
    .A1(_0474_),
    .S(net109),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1539_ (.A0(_0450_),
    .A1(_0454_),
    .S(net117),
    .X(_0480_));
 sky130_fd_sc_hd__inv_1 _1540_ (.A(net10),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_1 _1541_ (.A(net43),
    .Y(_0490_));
 sky130_fd_sc_hd__and2_0 _1542_ (.A(_0494_),
    .B(_0492_),
    .X(_0491_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1543_ (.A(_0494_),
    .SLEEP(_0492_),
    .X(_0495_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1544_ (.A(_0496_),
    .SLEEP(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__and2_0 _1545_ (.A(_0494_),
    .B(_0492_),
    .X(_0496_));
 sky130_fd_sc_hd__xor2_1 _1546_ (.A(_0494_),
    .B(_0492_),
    .X(_0500_));
 sky130_fd_sc_hd__and2_0 _1547_ (.A(_0500_),
    .B(_0457_),
    .X(_0497_));
 sky130_fd_sc_hd__xor2_1 _1548_ (.A(_0457_),
    .B(_0500_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _1549_ (.A0(net10),
    .A1(_0489_),
    .S(net126),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(net43),
    .A1(_0490_),
    .S(net123),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _1551_ (.A0(_0504_),
    .A1(net128),
    .S(net118),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(_0521_),
    .A1(_0515_),
    .S(net110),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1553_ (.A0(_0491_),
    .A1(_0495_),
    .S(net118),
    .X(_0521_));
 sky130_fd_sc_hd__inv_1 _1554_ (.A(net11),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_1 _1555_ (.A(net44),
    .Y(_0531_));
 sky130_fd_sc_hd__and2_0 _1556_ (.A(_0535_),
    .B(_0533_),
    .X(_0532_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1557_ (.A(_0535_),
    .SLEEP(_0533_),
    .X(_0536_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1558_ (.A(_0537_),
    .SLEEP(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__and2_0 _1559_ (.A(_0535_),
    .B(_0533_),
    .X(_0537_));
 sky130_fd_sc_hd__xor2_1 _1560_ (.A(_0535_),
    .B(_0533_),
    .X(_0541_));
 sky130_fd_sc_hd__and2_4 _1561_ (.A(_0498_),
    .B(_0541_),
    .X(_0538_));
 sky130_fd_sc_hd__xor2_1 _1562_ (.A(_0498_),
    .B(_0541_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _1563_ (.A0(net11),
    .A1(_0530_),
    .S(net127),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(net44),
    .A1(_0531_),
    .S(net123),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _1565_ (.A0(_0545_),
    .A1(net129),
    .S(net118),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _1566_ (.A0(_0562_),
    .A1(_0556_),
    .S(net110),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(_0532_),
    .A1(_0536_),
    .S(net118),
    .X(_0562_));
 sky130_fd_sc_hd__inv_1 _1568_ (.A(net12),
    .Y(_0571_));
 sky130_fd_sc_hd__inv_1 _1569_ (.A(net45),
    .Y(_0572_));
 sky130_fd_sc_hd__and2_0 _1570_ (.A(_0576_),
    .B(_0574_),
    .X(_0573_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1571_ (.A(_0576_),
    .SLEEP(_0574_),
    .X(_0577_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1572_ (.A(_0578_),
    .SLEEP(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__and2_0 _1573_ (.A(_0576_),
    .B(_0574_),
    .X(_0578_));
 sky130_fd_sc_hd__xor2_1 _1574_ (.A(_0576_),
    .B(_0574_),
    .X(_0582_));
 sky130_fd_sc_hd__and2_4 _1575_ (.A(_0088_),
    .B(_0582_),
    .X(_0579_));
 sky130_fd_sc_hd__xor2_1 _1576_ (.A(_0088_),
    .B(_0582_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _1577_ (.A0(net12),
    .A1(_0571_),
    .S(net124),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _1578_ (.A0(net45),
    .A1(_0572_),
    .S(net120),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _1579_ (.A0(_0586_),
    .A1(net130),
    .S(net111),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _1580_ (.A0(_0603_),
    .A1(_0597_),
    .S(net107),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1581_ (.A0(_0573_),
    .A1(_0577_),
    .S(net111),
    .X(_0603_));
 sky130_fd_sc_hd__inv_1 _1582_ (.A(net13),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_1 _1583_ (.A(net46),
    .Y(_0613_));
 sky130_fd_sc_hd__and2_0 _1584_ (.A(_0617_),
    .B(_0615_),
    .X(_0614_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1585_ (.A(_0617_),
    .SLEEP(_0615_),
    .X(_0618_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1586_ (.A(_0619_),
    .SLEEP(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__and2_0 _1587_ (.A(_0617_),
    .B(_0615_),
    .X(_0619_));
 sky130_fd_sc_hd__xor2_1 _1588_ (.A(_0617_),
    .B(_0615_),
    .X(_0623_));
 sky130_fd_sc_hd__and2_0 _1589_ (.A(_0539_),
    .B(_0623_),
    .X(_0620_));
 sky130_fd_sc_hd__xor2_1 _1590_ (.A(_0539_),
    .B(_0623_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _1591_ (.A0(net13),
    .A1(_0612_),
    .S(net127),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _1592_ (.A0(net46),
    .A1(_0613_),
    .S(net123),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _1593_ (.A0(_0627_),
    .A1(net131),
    .S(net118),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _1594_ (.A0(_0644_),
    .A1(_0638_),
    .S(net110),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1595_ (.A0(_0614_),
    .A1(_0618_),
    .S(net118),
    .X(_0644_));
 sky130_fd_sc_hd__inv_1 _1596_ (.A(net14),
    .Y(_0653_));
 sky130_fd_sc_hd__inv_1 _1597_ (.A(net47),
    .Y(_0654_));
 sky130_fd_sc_hd__and2_0 _1598_ (.A(_0658_),
    .B(_0656_),
    .X(_0655_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1599_ (.A(_0658_),
    .SLEEP(_0656_),
    .X(_0659_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1600_ (.A(_0660_),
    .SLEEP(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__and2_0 _1601_ (.A(_0658_),
    .B(_0656_),
    .X(_0660_));
 sky130_fd_sc_hd__xor2_1 _1602_ (.A(_0658_),
    .B(_0656_),
    .X(_0664_));
 sky130_fd_sc_hd__and2_4 _1603_ (.A(_0621_),
    .B(_0664_),
    .X(_0661_));
 sky130_fd_sc_hd__xor2_1 _1604_ (.A(_0621_),
    .B(_0664_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _1605_ (.A0(net14),
    .A1(_0653_),
    .S(net127),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(net47),
    .A1(_0654_),
    .S(net123),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(_0668_),
    .A1(net132),
    .S(net117),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(_0685_),
    .A1(_0679_),
    .S(net110),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1609_ (.A0(_0655_),
    .A1(_0659_),
    .S(net117),
    .X(_0685_));
 sky130_fd_sc_hd__inv_1 _1610_ (.A(net15),
    .Y(_0694_));
 sky130_fd_sc_hd__inv_1 _1611_ (.A(net48),
    .Y(_0695_));
 sky130_fd_sc_hd__and2_0 _1612_ (.A(_0699_),
    .B(_0697_),
    .X(_0696_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1613_ (.A(_0699_),
    .SLEEP(_0697_),
    .X(_0700_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1614_ (.A(_0701_),
    .SLEEP(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__and2_0 _1615_ (.A(_0699_),
    .B(_0697_),
    .X(_0701_));
 sky130_fd_sc_hd__xor2_1 _1616_ (.A(_0699_),
    .B(_0697_),
    .X(_0705_));
 sky130_fd_sc_hd__and2_0 _1617_ (.A(_0662_),
    .B(_0705_),
    .X(_0702_));
 sky130_fd_sc_hd__xor2_1 _1618_ (.A(net161),
    .B(_0705_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _1619_ (.A0(net15),
    .A1(_0694_),
    .S(net127),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _1620_ (.A0(net48),
    .A1(_0695_),
    .S(net123),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _1621_ (.A0(_0709_),
    .A1(net133),
    .S(net117),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _1622_ (.A0(_0726_),
    .A1(_0720_),
    .S(net110),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1623_ (.A0(_0696_),
    .A1(_0700_),
    .S(net117),
    .X(_0726_));
 sky130_fd_sc_hd__inv_1 _1624_ (.A(net16),
    .Y(_0735_));
 sky130_fd_sc_hd__inv_1 _1625_ (.A(net49),
    .Y(_0736_));
 sky130_fd_sc_hd__and2_0 _1626_ (.A(_0740_),
    .B(_0738_),
    .X(_0737_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1627_ (.A(_0740_),
    .SLEEP(_0738_),
    .X(_0741_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1628_ (.A(_0742_),
    .SLEEP(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__and2_0 _1629_ (.A(_0740_),
    .B(_0738_),
    .X(_0742_));
 sky130_fd_sc_hd__xor2_1 _1630_ (.A(_0740_),
    .B(_0738_),
    .X(_0746_));
 sky130_fd_sc_hd__and2_4 _1631_ (.A(_0703_),
    .B(_0746_),
    .X(_0743_));
 sky130_fd_sc_hd__xor2_1 _1632_ (.A(net163),
    .B(_0746_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _1633_ (.A0(net16),
    .A1(_0735_),
    .S(net125),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _1634_ (.A0(net49),
    .A1(_0736_),
    .S(net123),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _1635_ (.A0(_0750_),
    .A1(net134),
    .S(net117),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _1636_ (.A0(_0767_),
    .A1(_0761_),
    .S(net110),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1637_ (.A0(_0737_),
    .A1(_0741_),
    .S(net117),
    .X(_0767_));
 sky130_fd_sc_hd__inv_1 _1638_ (.A(net17),
    .Y(_0776_));
 sky130_fd_sc_hd__inv_1 _1639_ (.A(net50),
    .Y(_0777_));
 sky130_fd_sc_hd__and2_0 _1640_ (.A(_0781_),
    .B(_0779_),
    .X(_0778_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1641_ (.A(_0781_),
    .SLEEP(_0779_),
    .X(_0782_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1642_ (.A(_0783_),
    .SLEEP(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__and2_0 _1643_ (.A(_0781_),
    .B(_0779_),
    .X(_0783_));
 sky130_fd_sc_hd__xor2_1 _1644_ (.A(_0781_),
    .B(_0779_),
    .X(_0787_));
 sky130_fd_sc_hd__and2_0 _1645_ (.A(_0744_),
    .B(_0787_),
    .X(_0784_));
 sky130_fd_sc_hd__xor2_1 _1646_ (.A(net165),
    .B(_0787_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _1647_ (.A0(net17),
    .A1(_0776_),
    .S(net125),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _1648_ (.A0(net50),
    .A1(_0777_),
    .S(net159),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _1649_ (.A0(_0791_),
    .A1(net135),
    .S(net114),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _1650_ (.A0(_0808_),
    .A1(_0802_),
    .S(net107),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1651_ (.A0(_0778_),
    .A1(_0782_),
    .S(net114),
    .X(_0808_));
 sky130_fd_sc_hd__inv_1 _1652_ (.A(net18),
    .Y(_0817_));
 sky130_fd_sc_hd__inv_1 _1653_ (.A(net51),
    .Y(_0818_));
 sky130_fd_sc_hd__and2_0 _1654_ (.A(_0822_),
    .B(_0820_),
    .X(_0819_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1655_ (.A(_0822_),
    .SLEEP(_0820_),
    .X(_0823_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1656_ (.A(_0824_),
    .SLEEP(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__and2_0 _1657_ (.A(_0822_),
    .B(_0820_),
    .X(_0824_));
 sky130_fd_sc_hd__xor2_1 _1658_ (.A(_0822_),
    .B(_0820_),
    .X(_0828_));
 sky130_fd_sc_hd__and2_0 _1659_ (.A(_0785_),
    .B(_0828_),
    .X(_0825_));
 sky130_fd_sc_hd__xor2_1 _1660_ (.A(net168),
    .B(_0828_),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _1661_ (.A0(net18),
    .A1(_0817_),
    .S(net125),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _1662_ (.A0(net51),
    .A1(_0818_),
    .S(net159),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _1663_ (.A0(_0832_),
    .A1(net136),
    .S(net114),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _1664_ (.A0(_0849_),
    .A1(_0843_),
    .S(net108),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1665_ (.A0(_0819_),
    .A1(_0823_),
    .S(net114),
    .X(_0849_));
 sky130_fd_sc_hd__inv_1 _1666_ (.A(net19),
    .Y(_0858_));
 sky130_fd_sc_hd__inv_1 _1667_ (.A(net52),
    .Y(_0859_));
 sky130_fd_sc_hd__and2_0 _1668_ (.A(_0863_),
    .B(_0861_),
    .X(_0860_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1669_ (.A(_0863_),
    .SLEEP(_0861_),
    .X(_0864_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1670_ (.A(_0865_),
    .SLEEP(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__and2_0 _1671_ (.A(_0863_),
    .B(_0861_),
    .X(_0865_));
 sky130_fd_sc_hd__xor2_1 _1672_ (.A(_0863_),
    .B(_0861_),
    .X(_0869_));
 sky130_fd_sc_hd__and2_0 _1673_ (.A(_0826_),
    .B(_0869_),
    .X(_0866_));
 sky130_fd_sc_hd__xor2_1 _1674_ (.A(net169),
    .B(_0869_),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _1675_ (.A0(net19),
    .A1(_0858_),
    .S(net125),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _1676_ (.A0(net52),
    .A1(_0859_),
    .S(net121),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(_0873_),
    .A1(net137),
    .S(net114),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _1678_ (.A0(_0890_),
    .A1(_0884_),
    .S(net108),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1679_ (.A0(_0860_),
    .A1(_0864_),
    .S(net114),
    .X(_0890_));
 sky130_fd_sc_hd__inv_1 _1680_ (.A(net20),
    .Y(_0899_));
 sky130_fd_sc_hd__inv_1 _1681_ (.A(net53),
    .Y(_0900_));
 sky130_fd_sc_hd__and2_0 _1682_ (.A(_0904_),
    .B(_0902_),
    .X(_0901_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1683_ (.A(_0904_),
    .SLEEP(_0902_),
    .X(_0905_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1684_ (.A(_0906_),
    .SLEEP(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__and2_0 _1685_ (.A(_0904_),
    .B(_0902_),
    .X(_0906_));
 sky130_fd_sc_hd__xor2_1 _1686_ (.A(_0904_),
    .B(_0902_),
    .X(_0910_));
 sky130_fd_sc_hd__and2_0 _1687_ (.A(_0867_),
    .B(_0910_),
    .X(_0907_));
 sky130_fd_sc_hd__xor2_1 _1688_ (.A(net167),
    .B(_0910_),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _1689_ (.A0(net20),
    .A1(_0899_),
    .S(net125),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _1690_ (.A0(net53),
    .A1(_0900_),
    .S(net121),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _1691_ (.A0(_0914_),
    .A1(net138),
    .S(net113),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _1692_ (.A0(_0931_),
    .A1(_0925_),
    .S(net108),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1693_ (.A0(_0901_),
    .A1(_0905_),
    .S(net113),
    .X(_0931_));
 sky130_fd_sc_hd__inv_1 _1694_ (.A(net21),
    .Y(_0940_));
 sky130_fd_sc_hd__inv_1 _1695_ (.A(net54),
    .Y(_0941_));
 sky130_fd_sc_hd__and2_0 _1696_ (.A(_0945_),
    .B(_0943_),
    .X(_0942_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1697_ (.A(_0945_),
    .SLEEP(_0943_),
    .X(_0946_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1698_ (.A(_0947_),
    .SLEEP(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__and2_0 _1699_ (.A(_0945_),
    .B(_0943_),
    .X(_0947_));
 sky130_fd_sc_hd__xor2_1 _1700_ (.A(_0945_),
    .B(_0943_),
    .X(_0951_));
 sky130_fd_sc_hd__and2_0 _1701_ (.A(_0908_),
    .B(_0951_),
    .X(_0948_));
 sky130_fd_sc_hd__xor2_1 _1702_ (.A(net166),
    .B(_0951_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _1703_ (.A0(net21),
    .A1(_0940_),
    .S(net125),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(net54),
    .A1(_0941_),
    .S(net121),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(_0955_),
    .A1(net139),
    .S(net113),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _1706_ (.A0(_0972_),
    .A1(_0966_),
    .S(net108),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1707_ (.A0(_0942_),
    .A1(_0946_),
    .S(net113),
    .X(_0972_));
 sky130_fd_sc_hd__inv_1 _1708_ (.A(net22),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_1 _1709_ (.A(net55),
    .Y(_0982_));
 sky130_fd_sc_hd__and2_0 _1710_ (.A(_0986_),
    .B(_0984_),
    .X(_0983_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1711_ (.A(_0986_),
    .SLEEP(_0984_),
    .X(_0987_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1712_ (.A(_0988_),
    .SLEEP(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__and2_0 _1713_ (.A(_0986_),
    .B(_0984_),
    .X(_0988_));
 sky130_fd_sc_hd__xor2_1 _1714_ (.A(_0986_),
    .B(_0984_),
    .X(_0992_));
 sky130_fd_sc_hd__and2_0 _1715_ (.A(_0949_),
    .B(_0992_),
    .X(_0989_));
 sky130_fd_sc_hd__xor2_1 _1716_ (.A(net164),
    .B(_0992_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _1717_ (.A0(net22),
    .A1(_0981_),
    .S(net125),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _1718_ (.A0(net55),
    .A1(_0982_),
    .S(net121),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _1719_ (.A0(_0996_),
    .A1(net140),
    .S(net113),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _1720_ (.A0(_1013_),
    .A1(_1007_),
    .S(net108),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1721_ (.A0(_0983_),
    .A1(_0987_),
    .S(net113),
    .X(_1013_));
 sky130_fd_sc_hd__inv_1 _1722_ (.A(net23),
    .Y(_1022_));
 sky130_fd_sc_hd__inv_1 _1723_ (.A(net56),
    .Y(_1023_));
 sky130_fd_sc_hd__and2_0 _1724_ (.A(_1027_),
    .B(_1025_),
    .X(_1024_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1725_ (.A(_1027_),
    .SLEEP(_1025_),
    .X(_1028_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1726_ (.A(_1029_),
    .SLEEP(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__and2_0 _1727_ (.A(_1027_),
    .B(_1025_),
    .X(_1029_));
 sky130_fd_sc_hd__xor2_1 _1728_ (.A(_1027_),
    .B(_1025_),
    .X(_1033_));
 sky130_fd_sc_hd__and2_0 _1729_ (.A(_1033_),
    .B(_0580_),
    .X(_1030_));
 sky130_fd_sc_hd__xor2_1 _1730_ (.A(_0580_),
    .B(_1033_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _1731_ (.A0(net23),
    .A1(_1022_),
    .S(net124),
    .X(_1025_));
 sky130_fd_sc_hd__mux2_1 _1732_ (.A0(net56),
    .A1(_1023_),
    .S(net120),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_1 _1733_ (.A0(_1037_),
    .A1(net141),
    .S(net111),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _1734_ (.A0(_1054_),
    .A1(_1048_),
    .S(net107),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1735_ (.A0(_1024_),
    .A1(_1028_),
    .S(net111),
    .X(_1054_));
 sky130_fd_sc_hd__inv_1 _1736_ (.A(net24),
    .Y(_1063_));
 sky130_fd_sc_hd__inv_1 _1737_ (.A(net57),
    .Y(_1064_));
 sky130_fd_sc_hd__and2_0 _1738_ (.A(_1068_),
    .B(_1066_),
    .X(_1065_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1739_ (.A(_1068_),
    .SLEEP(_1066_),
    .X(_1069_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1740_ (.A(_1070_),
    .SLEEP(_1071_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_0 _1741_ (.A(_1068_),
    .B(_1066_),
    .X(_1070_));
 sky130_fd_sc_hd__xor2_1 _1742_ (.A(_1068_),
    .B(_1066_),
    .X(_1074_));
 sky130_fd_sc_hd__and2_4 _1743_ (.A(_0990_),
    .B(_1074_),
    .X(_1071_));
 sky130_fd_sc_hd__xor2_1 _1744_ (.A(net162),
    .B(_1074_),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_1 _1745_ (.A0(net24),
    .A1(_1063_),
    .S(net125),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _1746_ (.A0(net57),
    .A1(_1064_),
    .S(net121),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _1747_ (.A0(_1078_),
    .A1(net142),
    .S(net113),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_2 _1748_ (.A0(_1095_),
    .A1(_1089_),
    .S(net108),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1749_ (.A0(_1065_),
    .A1(_1069_),
    .S(net113),
    .X(_1095_));
 sky130_fd_sc_hd__inv_1 _1750_ (.A(net26),
    .Y(_1104_));
 sky130_fd_sc_hd__inv_1 _1751_ (.A(net59),
    .Y(_1105_));
 sky130_fd_sc_hd__and2_0 _1752_ (.A(_1109_),
    .B(_1107_),
    .X(_1106_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1753_ (.A(_1109_),
    .SLEEP(_1107_),
    .X(_1110_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1754_ (.A(_1111_),
    .SLEEP(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__and2_0 _1755_ (.A(_1109_),
    .B(_1107_),
    .X(_1111_));
 sky130_fd_sc_hd__xor2_1 _1756_ (.A(_1109_),
    .B(_1107_),
    .X(_1115_));
 sky130_fd_sc_hd__and2_4 _1757_ (.A(_1031_),
    .B(_1115_),
    .X(_1112_));
 sky130_fd_sc_hd__xor2_1 _1758_ (.A(_1031_),
    .B(_1115_),
    .X(_1119_));
 sky130_fd_sc_hd__mux2_1 _1759_ (.A0(net26),
    .A1(_1104_),
    .S(net124),
    .X(_1107_));
 sky130_fd_sc_hd__mux2_1 _1760_ (.A0(net59),
    .A1(_1105_),
    .S(net120),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _1761_ (.A0(_1119_),
    .A1(net143),
    .S(net111),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_1 _1762_ (.A0(_1136_),
    .A1(_1130_),
    .S(net107),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1763_ (.A0(_1106_),
    .A1(_1110_),
    .S(net111),
    .X(_1136_));
 sky130_fd_sc_hd__inv_1 _1764_ (.A(net27),
    .Y(_1145_));
 sky130_fd_sc_hd__inv_1 _1765_ (.A(net60),
    .Y(_1146_));
 sky130_fd_sc_hd__and2_0 _1766_ (.A(_1150_),
    .B(_1148_),
    .X(_1147_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1767_ (.A(_1150_),
    .SLEEP(_1148_),
    .X(_1151_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1768_ (.A(_1152_),
    .SLEEP(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__and2_0 _1769_ (.A(_1150_),
    .B(_1148_),
    .X(_1152_));
 sky130_fd_sc_hd__xor2_1 _1770_ (.A(_1150_),
    .B(_1148_),
    .X(_1156_));
 sky130_fd_sc_hd__and2_4 _1771_ (.A(_1113_),
    .B(_1156_),
    .X(_1153_));
 sky130_fd_sc_hd__xor2_1 _1772_ (.A(_1113_),
    .B(_1156_),
    .X(_1160_));
 sky130_fd_sc_hd__mux2_1 _1773_ (.A0(net27),
    .A1(_1145_),
    .S(net124),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _1774_ (.A0(net60),
    .A1(_1146_),
    .S(net120),
    .X(_1150_));
 sky130_fd_sc_hd__mux2_1 _1775_ (.A0(_1160_),
    .A1(net144),
    .S(net111),
    .X(_1171_));
 sky130_fd_sc_hd__mux2_1 _1776_ (.A0(_1177_),
    .A1(_1171_),
    .S(net107),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1777_ (.A0(_1147_),
    .A1(_1151_),
    .S(net111),
    .X(_1177_));
 sky130_fd_sc_hd__inv_1 _1778_ (.A(net28),
    .Y(_1186_));
 sky130_fd_sc_hd__inv_1 _1779_ (.A(net61),
    .Y(_1187_));
 sky130_fd_sc_hd__and2_0 _1780_ (.A(_1191_),
    .B(_1189_),
    .X(_1188_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1781_ (.A(_1191_),
    .SLEEP(_1189_),
    .X(_1192_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1782_ (.A(_1193_),
    .SLEEP(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__and2_0 _1783_ (.A(_1191_),
    .B(_1189_),
    .X(_1193_));
 sky130_fd_sc_hd__xor2_1 _1784_ (.A(_1191_),
    .B(_1189_),
    .X(_1197_));
 sky130_fd_sc_hd__and2_4 _1785_ (.A(_1154_),
    .B(_1197_),
    .X(_1194_));
 sky130_fd_sc_hd__xor2_1 _1786_ (.A(_1154_),
    .B(_1197_),
    .X(_1201_));
 sky130_fd_sc_hd__mux2_1 _1787_ (.A0(net28),
    .A1(_1186_),
    .S(net160),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _1788_ (.A0(net61),
    .A1(_1187_),
    .S(net159),
    .X(_1191_));
 sky130_fd_sc_hd__mux2_1 _1789_ (.A0(_1201_),
    .A1(net145),
    .S(net112),
    .X(_1212_));
 sky130_fd_sc_hd__mux2_1 _1790_ (.A0(_1218_),
    .A1(_1212_),
    .S(net107),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1791_ (.A0(_1188_),
    .A1(_1192_),
    .S(net112),
    .X(_1218_));
 sky130_fd_sc_hd__inv_1 _1792_ (.A(net29),
    .Y(_1227_));
 sky130_fd_sc_hd__inv_1 _1793_ (.A(net62),
    .Y(_1228_));
 sky130_fd_sc_hd__and2_0 _1794_ (.A(_1232_),
    .B(_1230_),
    .X(_1229_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1795_ (.A(_1232_),
    .SLEEP(_1230_),
    .X(_1233_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1796_ (.A(_1234_),
    .SLEEP(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__and2_0 _1797_ (.A(_1232_),
    .B(_1230_),
    .X(_1234_));
 sky130_fd_sc_hd__xor2_1 _1798_ (.A(_1232_),
    .B(_1230_),
    .X(_1238_));
 sky130_fd_sc_hd__and2_4 _1799_ (.A(_1195_),
    .B(_1238_),
    .X(_1235_));
 sky130_fd_sc_hd__xor2_1 _1800_ (.A(_1195_),
    .B(_1238_),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _1801_ (.A0(net29),
    .A1(_1227_),
    .S(net160),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _1802_ (.A0(net62),
    .A1(_1228_),
    .S(net159),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _1803_ (.A0(_1242_),
    .A1(net146),
    .S(net112),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_1 _1804_ (.A0(_1259_),
    .A1(_1253_),
    .S(net107),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(_1229_),
    .A1(_1233_),
    .S(net112),
    .X(_1259_));
 sky130_fd_sc_hd__inv_1 _1806_ (.A(net30),
    .Y(_1268_));
 sky130_fd_sc_hd__inv_1 _1807_ (.A(net63),
    .Y(_1269_));
 sky130_fd_sc_hd__and2_0 _1808_ (.A(_1273_),
    .B(_1271_),
    .X(_1270_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1809_ (.A(_1273_),
    .SLEEP(_1271_),
    .X(_1274_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1810_ (.A(_1275_),
    .SLEEP(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__and2_0 _1811_ (.A(_1273_),
    .B(_1271_),
    .X(_1275_));
 sky130_fd_sc_hd__xor2_1 _1812_ (.A(_1273_),
    .B(_1271_),
    .X(_1279_));
 sky130_fd_sc_hd__and2_0 _1813_ (.A(_1236_),
    .B(_1279_),
    .X(_1276_));
 sky130_fd_sc_hd__xor2_1 _1814_ (.A(_1236_),
    .B(_1279_),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _1815_ (.A0(net30),
    .A1(_1268_),
    .S(net160),
    .X(_1271_));
 sky130_fd_sc_hd__mux2_1 _1816_ (.A0(net63),
    .A1(_1269_),
    .S(net121),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _1817_ (.A0(_1283_),
    .A1(net147),
    .S(net112),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _1818_ (.A0(_1300_),
    .A1(_1294_),
    .S(net107),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1819_ (.A0(_1270_),
    .A1(_1274_),
    .S(net112),
    .X(_1300_));
 sky130_fd_sc_hd__inv_1 _1820_ (.A(net31),
    .Y(_1309_));
 sky130_fd_sc_hd__inv_1 _1821_ (.A(net64),
    .Y(_1310_));
 sky130_fd_sc_hd__and2_0 _1822_ (.A(_1314_),
    .B(_1312_),
    .X(_1311_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1823_ (.A(_1314_),
    .SLEEP(_1312_),
    .X(_1315_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1824_ (.A(_1316_),
    .SLEEP(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__and2_0 _1825_ (.A(_1314_),
    .B(_1312_),
    .X(_1316_));
 sky130_fd_sc_hd__xor2_1 _1826_ (.A(_1314_),
    .B(_1312_),
    .X(_1320_));
 sky130_fd_sc_hd__and2_4 _1827_ (.A(_1277_),
    .B(_1320_),
    .X(_1317_));
 sky130_fd_sc_hd__xor2_1 _1828_ (.A(_1277_),
    .B(_1320_),
    .X(_1324_));
 sky130_fd_sc_hd__mux2_1 _1829_ (.A0(net31),
    .A1(_1309_),
    .S(net126),
    .X(_1312_));
 sky130_fd_sc_hd__mux2_1 _1830_ (.A0(net64),
    .A1(_1310_),
    .S(net122),
    .X(_1314_));
 sky130_fd_sc_hd__mux2_1 _1831_ (.A0(_1324_),
    .A1(net148),
    .S(net115),
    .X(_1335_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(_1341_),
    .A1(_1335_),
    .S(net109),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1833_ (.A0(_1311_),
    .A1(_1315_),
    .S(net115),
    .X(_1341_));
 sky130_fd_sc_hd__inv_1 _1834_ (.A(net32),
    .Y(_1350_));
 sky130_fd_sc_hd__inv_1 _1835_ (.A(net65),
    .Y(_1351_));
 sky130_fd_sc_hd__and2_0 _1836_ (.A(_1355_),
    .B(_1353_),
    .X(_1352_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1837_ (.A(_1355_),
    .SLEEP(_1353_),
    .X(_1356_));
 sky130_fd_sc_hd__lpflow_inputiso1p_1 _1838_ (.A(_1357_),
    .SLEEP(_1358_),
    .X(_0178_));
 sky130_fd_sc_hd__and2_0 _1839_ (.A(_1355_),
    .B(_1353_),
    .X(_1357_));
 sky130_fd_sc_hd__xor2_1 _1840_ (.A(_1355_),
    .B(_1353_),
    .X(_1361_));
 sky130_fd_sc_hd__and2_4 _1841_ (.A(_1318_),
    .B(_1361_),
    .X(_1358_));
 sky130_fd_sc_hd__xor2_1 _1842_ (.A(_1318_),
    .B(_1361_),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_1 _1843_ (.A0(net32),
    .A1(_1350_),
    .S(net160),
    .X(_1353_));
 sky130_fd_sc_hd__mux2_1 _1844_ (.A0(net65),
    .A1(_1351_),
    .S(net122),
    .X(_1355_));
 sky130_fd_sc_hd__mux2_1 _1845_ (.A0(_1365_),
    .A1(net149),
    .S(net115),
    .X(_1376_));
 sky130_fd_sc_hd__mux2_1 _1846_ (.A0(_1382_),
    .A1(_1376_),
    .S(net109),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1847_ (.A0(_1352_),
    .A1(_1356_),
    .S(net115),
    .X(_1382_));
 sky130_fd_sc_hd__conb_1 _1565__129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 _1579__130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 _1593__131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 _1607__132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 _1621__133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 _1635__134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 _1649__135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 _1663__136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 _1677__137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 _1691__138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 _1705__139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 _1719__140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 _1733__141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 _1747__142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 _1761__143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 _1775__144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 _1789__145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 _1803__146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 _1817__147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 _1831__148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 _1845__149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 _1425__150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 _1439__151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 _1453__152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 _1467__153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 _1481__154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 _1495__155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 _1509__156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 _1523__157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 _1537__158 (.LO(net158));
 sky130_fd_sc_hd__clkbuf_16 clone1 (.A(net66),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _1910_ (.A(_0043_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _1911_ (.A(_0054_),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _1912_ (.A(_0065_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _1913_ (.A(_0068_),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _1914_ (.A(_0069_),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _1915_ (.A(_0070_),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _1916_ (.A(_0071_),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _1917_ (.A(_0072_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _1918_ (.A(_0073_),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _1919_ (.A(_0074_),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _1920_ (.A(_0044_),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _1921_ (.A(_0045_),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _1922_ (.A(_0046_),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _1923_ (.A(_0047_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _1924_ (.A(_0048_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _1925_ (.A(_0049_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _1926_ (.A(_0050_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _1927_ (.A(_0051_),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _1928_ (.A(_0052_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _1929_ (.A(_0053_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _1930_ (.A(_0055_),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _1931_ (.A(_0056_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _1932_ (.A(_0057_),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _1933_ (.A(_0058_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _1934_ (.A(_0059_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _1935_ (.A(_0060_),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _1936_ (.A(_0061_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _1937_ (.A(_0062_),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _1938_ (.A(_0063_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _1939_ (.A(_0064_),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _1940_ (.A(_0066_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _1941_ (.A(_0067_),
    .X(net96));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_241 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(ainv),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(b[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(b[10]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(b[11]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(b[12]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(b[13]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(b[14]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(b[15]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(b[16]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(b[17]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(b[18]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(b[19]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(b[1]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(b[20]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(b[21]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(b[22]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(b[23]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(b[24]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(b[25]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(b[26]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(b[27]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(b[28]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(b[29]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(b[2]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(b[30]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(b[31]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(b[3]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b[4]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b[5]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b[6]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(b[7]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(b[8]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(b[9]),
    .X(net65));
 sky130_fd_sc_hd__buf_6 input66 (.A(binv),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(cin),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(select[0]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(select[1]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(cout));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(overflow));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(result[0]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(result[10]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(result[11]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(result[12]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(result[13]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(result[14]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(result[15]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(result[16]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(result[17]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(result[18]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(result[19]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(result[1]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(result[20]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(result[21]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(result[22]));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net87),
    .X(result[23]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(result[24]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(result[25]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(result[26]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(result[27]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(result[28]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(result[29]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(result[2]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(result[30]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(result[31]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(result[3]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(result[4]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(result[5]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(result[6]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(result[7]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(result[8]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(result[9]));
 sky130_fd_sc_hd__buf_4 output104 (.A(net104),
    .X(zero));
 sky130_fd_sc_hd__clkbuf_1 wire105 (.A(_0040_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 wire106 (.A(_0035_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(net69),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 fanout108 (.A(net69),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 fanout109 (.A(net69),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(net69),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net119),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(net119),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net119),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 fanout114 (.A(net119),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net119),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 fanout116 (.A(net119),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(net119),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(net68),
    .X(net119));
 sky130_fd_sc_hd__buf_8 fanout120 (.A(net66),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net66),
    .X(net121));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net66),
    .X(net122));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(net66),
    .X(net123));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(net127),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(net127),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_8 fanout127 (.A(net33),
    .X(net127));
 sky130_fd_sc_hd__conb_1 _1551__128 (.LO(net128));
 sky130_fd_sc_hd__clkbuf_16 clone2 (.A(net127),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(_0662_),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(_0990_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_0703_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(_0949_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(_0744_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(_0908_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(_0867_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(_0785_),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(_0826_),
    .X(net169));
endmodule
