magic
tech sky130A
magscale 1 2
timestamp 1743983954
<< nwell >>
rect 1066 2159 22394 23430
<< obsli1 >>
rect 1104 2159 22356 23409
<< obsm1 >>
rect 842 2128 22356 23440
<< metal2 >>
rect 4526 24812 4582 25612
rect 5170 24812 5226 25612
rect 6458 24812 6514 25612
rect 7102 24812 7158 25612
rect 7746 24812 7802 25612
rect 8390 24812 8446 25612
rect 9034 24812 9090 25612
rect 9678 24812 9734 25612
rect 10322 24812 10378 25612
rect 10966 24812 11022 25612
rect 11610 24812 11666 25612
rect 12254 24812 12310 25612
rect 12898 24812 12954 25612
rect 13542 24812 13598 25612
rect 14186 24812 14242 25612
rect 14830 24812 14886 25612
rect 15474 24812 15530 25612
rect 16118 24812 16174 25612
rect 16762 24812 16818 25612
rect 17406 24812 17462 25612
rect 18050 24812 18106 25612
rect 18694 24812 18750 25612
rect 19338 24812 19394 25612
rect 18 0 74 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
<< obsm2 >>
rect 846 24756 4470 24970
rect 4638 24756 5114 24970
rect 5282 24756 6402 24970
rect 6570 24756 7046 24970
rect 7214 24756 7690 24970
rect 7858 24756 8334 24970
rect 8502 24756 8978 24970
rect 9146 24756 9622 24970
rect 9790 24756 10266 24970
rect 10434 24756 10910 24970
rect 11078 24756 11554 24970
rect 11722 24756 12198 24970
rect 12366 24756 12842 24970
rect 13010 24756 13486 24970
rect 13654 24756 14130 24970
rect 14298 24756 14774 24970
rect 14942 24756 15418 24970
rect 15586 24756 16062 24970
rect 16230 24756 16706 24970
rect 16874 24756 17350 24970
rect 17518 24756 17994 24970
rect 18162 24756 18638 24970
rect 18806 24756 19282 24970
rect 19450 24756 22062 24970
rect 846 856 22062 24756
rect 846 734 3182 856
rect 3350 734 3826 856
rect 3994 734 4470 856
rect 4638 734 5114 856
rect 5282 734 5758 856
rect 5926 734 6402 856
rect 6570 734 7046 856
rect 7214 734 7690 856
rect 7858 734 8334 856
rect 8502 734 8978 856
rect 9146 734 9622 856
rect 9790 734 10266 856
rect 10434 734 10910 856
rect 11078 734 11554 856
rect 11722 734 12198 856
rect 12366 734 12842 856
rect 13010 734 13486 856
rect 13654 734 14130 856
rect 14298 734 14774 856
rect 14942 734 15418 856
rect 15586 734 16062 856
rect 16230 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17994 856
rect 18162 734 18638 856
rect 18806 734 19282 856
rect 19450 734 19926 856
rect 20094 734 22062 856
<< metal3 >>
rect 0 22448 800 22568
rect 0 21768 800 21888
rect 0 21088 800 21208
rect 0 20408 800 20528
rect 22668 20408 23468 20528
rect 0 19728 800 19848
rect 22668 19728 23468 19848
rect 0 19048 800 19168
rect 22668 19048 23468 19168
rect 0 18368 800 18488
rect 22668 18368 23468 18488
rect 0 17688 800 17808
rect 22668 17688 23468 17808
rect 0 17008 800 17128
rect 22668 17008 23468 17128
rect 0 16328 800 16448
rect 22668 16328 23468 16448
rect 0 15648 800 15768
rect 22668 15648 23468 15768
rect 0 14968 800 15088
rect 22668 14968 23468 15088
rect 0 14288 800 14408
rect 22668 14288 23468 14408
rect 0 13608 800 13728
rect 22668 13608 23468 13728
rect 0 12928 800 13048
rect 22668 12928 23468 13048
rect 0 12248 800 12368
rect 22668 12248 23468 12368
rect 0 11568 800 11688
rect 22668 11568 23468 11688
rect 0 10888 800 11008
rect 22668 10888 23468 11008
rect 0 10208 800 10328
rect 22668 10208 23468 10328
rect 0 9528 800 9648
rect 22668 9528 23468 9648
rect 0 8848 800 8968
rect 22668 8848 23468 8968
rect 0 8168 800 8288
rect 22668 8168 23468 8288
rect 0 7488 800 7608
rect 22668 7488 23468 7608
rect 0 6808 800 6928
rect 22668 6808 23468 6928
rect 0 6128 800 6248
rect 22668 6128 23468 6248
rect 0 5448 800 5568
rect 22668 5448 23468 5568
rect 0 4768 800 4888
rect 22668 4768 23468 4888
rect 0 4088 800 4208
rect 22668 4088 23468 4208
rect 0 3408 800 3528
<< obsm3 >>
rect 798 22648 22668 23425
rect 880 22368 22668 22648
rect 798 21968 22668 22368
rect 880 21688 22668 21968
rect 798 21288 22668 21688
rect 880 21008 22668 21288
rect 798 20608 22668 21008
rect 880 20328 22588 20608
rect 798 19928 22668 20328
rect 880 19648 22588 19928
rect 798 19248 22668 19648
rect 880 18968 22588 19248
rect 798 18568 22668 18968
rect 880 18288 22588 18568
rect 798 17888 22668 18288
rect 880 17608 22588 17888
rect 798 17208 22668 17608
rect 880 16928 22588 17208
rect 798 16528 22668 16928
rect 880 16248 22588 16528
rect 798 15848 22668 16248
rect 880 15568 22588 15848
rect 798 15168 22668 15568
rect 880 14888 22588 15168
rect 798 14488 22668 14888
rect 880 14208 22588 14488
rect 798 13808 22668 14208
rect 880 13528 22588 13808
rect 798 13128 22668 13528
rect 880 12848 22588 13128
rect 798 12448 22668 12848
rect 880 12168 22588 12448
rect 798 11768 22668 12168
rect 880 11488 22588 11768
rect 798 11088 22668 11488
rect 880 10808 22588 11088
rect 798 10408 22668 10808
rect 880 10128 22588 10408
rect 798 9728 22668 10128
rect 880 9448 22588 9728
rect 798 9048 22668 9448
rect 880 8768 22588 9048
rect 798 8368 22668 8768
rect 880 8088 22588 8368
rect 798 7688 22668 8088
rect 880 7408 22588 7688
rect 798 7008 22668 7408
rect 880 6728 22588 7008
rect 798 6328 22668 6728
rect 880 6048 22588 6328
rect 798 5648 22668 6048
rect 880 5368 22588 5648
rect 798 4968 22668 5368
rect 880 4688 22588 4968
rect 798 4288 22668 4688
rect 880 4008 22588 4288
rect 798 3608 22668 4008
rect 880 3328 22668 3608
rect 798 2143 22668 3328
<< metal4 >>
rect 3600 2128 3920 23440
rect 4260 2128 4580 23440
rect 8913 2128 9233 23440
rect 9573 2128 9893 23440
rect 14226 2128 14546 23440
rect 14886 2128 15206 23440
rect 19539 2128 19859 23440
rect 20199 2128 20519 23440
<< metal5 >>
rect 1056 21240 22404 21560
rect 1056 20580 22404 20900
rect 1056 15936 22404 16256
rect 1056 15276 22404 15596
rect 1056 10632 22404 10952
rect 1056 9972 22404 10292
rect 1056 5328 22404 5648
rect 1056 4668 22404 4988
<< labels >>
rlabel metal4 s 4260 2128 4580 23440 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 9573 2128 9893 23440 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 14886 2128 15206 23440 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 20199 2128 20519 23440 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5328 22404 5648 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 10632 22404 10952 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 15936 22404 16256 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 21240 22404 21560 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3600 2128 3920 23440 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8913 2128 9233 23440 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 14226 2128 14546 23440 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19539 2128 19859 23440 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4668 22404 4988 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 9972 22404 10292 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 15276 22404 15596 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 20580 22404 20900 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 3238 0 3294 800 6 a[0]
port 3 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 a[10]
port 4 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 a[11]
port 5 nsew signal input
rlabel metal2 s 5170 24812 5226 25612 6 a[12]
port 6 nsew signal input
rlabel metal2 s 8390 24812 8446 25612 6 a[13]
port 7 nsew signal input
rlabel metal2 s 9034 24812 9090 25612 6 a[14]
port 8 nsew signal input
rlabel metal2 s 10966 24812 11022 25612 6 a[15]
port 9 nsew signal input
rlabel metal2 s 15474 24812 15530 25612 6 a[16]
port 10 nsew signal input
rlabel metal2 s 13542 24812 13598 25612 6 a[17]
port 11 nsew signal input
rlabel metal2 s 18694 24812 18750 25612 6 a[18]
port 12 nsew signal input
rlabel metal3 s 22668 20408 23468 20528 6 a[19]
port 13 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 a[1]
port 14 nsew signal input
rlabel metal3 s 22668 19728 23468 19848 6 a[20]
port 15 nsew signal input
rlabel metal3 s 22668 15648 23468 15768 6 a[21]
port 16 nsew signal input
rlabel metal3 s 22668 19048 23468 19168 6 a[22]
port 17 nsew signal input
rlabel metal3 s 22668 12248 23468 12368 6 a[23]
port 18 nsew signal input
rlabel metal3 s 22668 11568 23468 11688 6 a[24]
port 19 nsew signal input
rlabel metal3 s 22668 14288 23468 14408 6 a[25]
port 20 nsew signal input
rlabel metal3 s 22668 4768 23468 4888 6 a[26]
port 21 nsew signal input
rlabel metal3 s 22668 5448 23468 5568 6 a[27]
port 22 nsew signal input
rlabel metal3 s 22668 4088 23468 4208 6 a[28]
port 23 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 a[29]
port 24 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 a[2]
port 25 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 a[30]
port 26 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 a[31]
port 27 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 a[3]
port 28 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 a[4]
port 29 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 a[5]
port 30 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 a[6]
port 31 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 a[7]
port 32 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 a[8]
port 33 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 a[9]
port 34 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 ainv
port 35 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 b[0]
port 36 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 b[10]
port 37 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 b[11]
port 38 nsew signal input
rlabel metal2 s 4526 24812 4582 25612 6 b[12]
port 39 nsew signal input
rlabel metal2 s 6458 24812 6514 25612 6 b[13]
port 40 nsew signal input
rlabel metal2 s 9678 24812 9734 25612 6 b[14]
port 41 nsew signal input
rlabel metal2 s 10322 24812 10378 25612 6 b[15]
port 42 nsew signal input
rlabel metal2 s 14830 24812 14886 25612 6 b[16]
port 43 nsew signal input
rlabel metal2 s 12898 24812 12954 25612 6 b[17]
port 44 nsew signal input
rlabel metal2 s 17406 24812 17462 25612 6 b[18]
port 45 nsew signal input
rlabel metal2 s 19338 24812 19394 25612 6 b[19]
port 46 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 b[1]
port 47 nsew signal input
rlabel metal3 s 22668 18368 23468 18488 6 b[20]
port 48 nsew signal input
rlabel metal3 s 22668 14968 23468 15088 6 b[21]
port 49 nsew signal input
rlabel metal3 s 22668 16328 23468 16448 6 b[22]
port 50 nsew signal input
rlabel metal3 s 22668 13608 23468 13728 6 b[23]
port 51 nsew signal input
rlabel metal3 s 22668 10888 23468 11008 6 b[24]
port 52 nsew signal input
rlabel metal3 s 22668 12928 23468 13048 6 b[25]
port 53 nsew signal input
rlabel metal3 s 22668 10208 23468 10328 6 b[26]
port 54 nsew signal input
rlabel metal3 s 22668 6808 23468 6928 6 b[27]
port 55 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 b[28]
port 56 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 b[29]
port 57 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 b[2]
port 58 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 b[30]
port 59 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 b[31]
port 60 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 b[3]
port 61 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 b[4]
port 62 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 b[5]
port 63 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 b[6]
port 64 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 b[7]
port 65 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 b[8]
port 66 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 b[9]
port 67 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 binv
port 68 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 cin
port 69 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 cout
port 70 nsew signal output
rlabel metal2 s 18 0 74 800 6 fake_clk
port 71 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 overflow
port 72 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 result[0]
port 73 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 result[10]
port 74 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 result[11]
port 75 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 result[12]
port 76 nsew signal output
rlabel metal2 s 7102 24812 7158 25612 6 result[13]
port 77 nsew signal output
rlabel metal2 s 7746 24812 7802 25612 6 result[14]
port 78 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 result[15]
port 79 nsew signal output
rlabel metal2 s 18050 24812 18106 25612 6 result[16]
port 80 nsew signal output
rlabel metal2 s 12254 24812 12310 25612 6 result[17]
port 81 nsew signal output
rlabel metal2 s 14186 24812 14242 25612 6 result[18]
port 82 nsew signal output
rlabel metal2 s 16118 24812 16174 25612 6 result[19]
port 83 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 result[1]
port 84 nsew signal output
rlabel metal2 s 16762 24812 16818 25612 6 result[20]
port 85 nsew signal output
rlabel metal3 s 22668 17688 23468 17808 6 result[21]
port 86 nsew signal output
rlabel metal3 s 22668 17008 23468 17128 6 result[22]
port 87 nsew signal output
rlabel metal2 s 11610 24812 11666 25612 6 result[23]
port 88 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 result[24]
port 89 nsew signal output
rlabel metal3 s 22668 6128 23468 6248 6 result[25]
port 90 nsew signal output
rlabel metal3 s 22668 9528 23468 9648 6 result[26]
port 91 nsew signal output
rlabel metal3 s 22668 7488 23468 7608 6 result[27]
port 92 nsew signal output
rlabel metal3 s 22668 8168 23468 8288 6 result[28]
port 93 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 result[29]
port 94 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 result[2]
port 95 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 result[30]
port 96 nsew signal output
rlabel metal3 s 22668 8848 23468 8968 6 result[31]
port 97 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 result[3]
port 98 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 result[4]
port 99 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 result[5]
port 100 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 result[6]
port 101 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 result[7]
port 102 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 result[8]
port 103 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 result[9]
port 104 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 select[0]
port 105 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 select[1]
port 106 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 zero
port 107 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 23468 25612
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1477886
string GDS_FILE /home/prajuval/Desktop/OpenLane/openlane/n_bit_alu/runs/run_8/results/signoff/n_bit_alu.magic.gds
string GDS_START 174250
<< end >>

