* NGSPICE file created from n_bit_alu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_0 abstract view
.subckt sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__lpflow_inputiso1p_1 abstract view
.subckt sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

.subckt n_bit_alu VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16] a[17] a[18]
+ a[19] a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29] a[2] a[30]
+ a[31] a[3] a[4] a[5] a[6] a[7] a[8] a[9] ainv b[0] b[10] b[11] b[12] b[13] b[14]
+ b[15] b[16] b[17] b[18] b[19] b[1] b[20] b[21] b[22] b[23] b[24] b[25] b[26] b[27]
+ b[28] b[29] b[2] b[30] b[31] b[3] b[4] b[5] b[6] b[7] b[8] b[9] binv cin cout fake_clk
+ overflow result[0] result[10] result[11] result[12] result[13] result[14] result[15]
+ result[16] result[17] result[18] result[19] result[1] result[20] result[21] result[22]
+ result[23] result[24] result[25] result[26] result[27] result[28] result[29] result[2]
+ result[30] result[31] result[3] result[4] result[5] result[6] result[7] result[8]
+ result[9] select[0] select[1] zero
XTAP_TAPCELL_ROW_9_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1606_ net47 _0654_ net66 VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1537_ _0463_ net135 net68 VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
X_1399_ net70 _0030_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__xor2_1
X_1468_ _0275_ _0269_ net69 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1940_ _0066_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1785_ _1154_ _1197_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__and2_0
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1923_ _0047_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1570_ _0576_ _0574_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__and2_0
XFILLER_0_21_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1768_ _1152_ _1153_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1837_ _1355_ _1353_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1699_ _0945_ _0943_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__and2_0
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput75 net75 VGND VGND VPWR VPWR result[12] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_33_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput86 net86 VGND VGND VPWR VPWR result[22] sky130_fd_sc_hd__buf_1
Xoutput97 net97 VGND VGND VPWR VPWR result[3] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_26_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1622_ _0726_ _0720_ net69 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_1
X_1553_ _0491_ _0495_ net68 VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__mux2_1
X_1484_ net6 VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__inv_1
XFILLER_0_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1536_ net42 _0449_ net66 VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux2_1
X_1605_ net14 _0653_ net33 VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__mux2_1
X_1398_ _0036_ _0041_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__nor2_1
X_1467_ _0258_ net130 net68 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1519_ _0375_ _0418_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and2_0
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1922_ _0046_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
X_1784_ _1191_ _1189_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1698_ _0947_ _0948_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1767_ _1150_ _1148_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_12_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1836_ _1355_ _1353_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__and2_0
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput87 net87 VGND VGND VPWR VPWR result[23] sky130_fd_sc_hd__buf_1
Xoutput76 net76 VGND VGND VPWR VPWR result[13] sky130_fd_sc_hd__buf_1
Xoutput98 net98 VGND VGND VPWR VPWR result[4] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_26_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1621_ _0709_ net110 net68 VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux2_1
X_1552_ _0521_ _0515_ net69 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux2_1
X_1483_ _0286_ _0290_ net68 VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
X_1803__123 VGND VGND VPWR VPWR _1803__123/HI net123 sky130_fd_sc_hd__conb_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1819_ _1270_ _1274_ net68 VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1535_ net9 _0448_ net33 VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1604_ _0621_ _0664_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__xor2_1
X_1466_ net37 _0244_ net66 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
X_1397_ _0037_ _0038_ _0039_ _0040_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__nand4_1
XFILLER_0_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1518_ _0412_ _0410_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__xor2_1
X_1449_ _0170_ _0213_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__and2_0
XFILLER_0_37_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1551__105 VGND VGND VPWR VPWR _1551__105/HI net105 sky130_fd_sc_hd__conb_1
X_1921_ _0045_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
X_1783_ _1191_ _1189_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__and2_0
XFILLER_0_21_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1691__115 VGND VGND VPWR VPWR _1691__115/HI net115 sky130_fd_sc_hd__conb_1
X_1835_ net65 VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__inv_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1697_ _0945_ _0943_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1766_ _1150_ _1148_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__and2_0
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput77 net77 VGND VGND VPWR VPWR result[14] sky130_fd_sc_hd__buf_1
Xoutput88 net88 VGND VGND VPWR VPWR result[24] sky130_fd_sc_hd__buf_1
Xoutput99 net99 VGND VGND VPWR VPWR result[5] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_26_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1551_ _0504_ net105 net68 VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__mux2_1
X_1620_ net48 _0695_ net66 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__mux2_1
X_1482_ _0316_ _0310_ net69 VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1818_ _1300_ _1294_ net69 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1749_ _1065_ _1069_ net68 VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__mux2_1
X_1465_ net4 _0243_ net33 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1603_ _0621_ _0664_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__and2_0
X_1534_ _0416_ _0459_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__xor2_1
X_1396_ _0074_ _0044_ _0046_ _0049_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_5_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1517_ _0412_ _0410_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__and2_0
X_1448_ _0207_ _0205_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1920_ _0044_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
X_1782_ _1193_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1765_ net60 VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__inv_1
X_1834_ net32 VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__inv_1
X_1696_ _0945_ _0943_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__and2_0
XFILLER_0_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput78 net78 VGND VGND VPWR VPWR result[15] sky130_fd_sc_hd__buf_1
Xoutput89 net89 VGND VGND VPWR VPWR result[25] sky130_fd_sc_hd__buf_1
XFILLER_0_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ net43 _0490_ net66 VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux2_1
X_1481_ _0299_ net131 net68 VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1748_ _1095_ _1089_ net69 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__mux2_1
X_1817_ _1283_ net124 net68 VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__mux2_1
X_1679_ _0860_ _0864_ net68 VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_37_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1602_ _0658_ _0656_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1533_ _0416_ _0459_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__and2_0
XFILLER_0_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1395_ _0043_ _0068_ _0070_ _0071_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__nor4_1
X_1464_ _0211_ _0254_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_20_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1516_ _0414_ _0415_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1447_ _0207_ _0205_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__and2_0
XFILLER_0_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1719__117 VGND VGND VPWR VPWR _1719__117/HI net117 sky130_fd_sc_hd__conb_1
X_1781_ _1191_ _1189_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_27_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1764_ net27 VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__inv_1
XFILLER_0_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1833_ _1311_ _1315_ net68 VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__mux2_1
X_1695_ net54 VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__inv_1
XFILLER_0_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput79 net79 VGND VGND VPWR VPWR result[16] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1480_ net38 _0285_ net66 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1747_ _1078_ net119 net68 VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__mux2_1
X_1678_ _0890_ _0884_ net69 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux2_1
X_1816_ net63 _1269_ net66 VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1532_ _0453_ _0451_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1601_ _0658_ _0656_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__and2_0
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1394_ _0059_ _0062_ _0064_ _0066_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__nor4_1
X_1463_ _0211_ _0254_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__and2_0
XTAP_TAPCELL_ROW_37_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1515_ _0412_ _0410_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1446_ _0209_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1429_ net35 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_41_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1780_ _1191_ _1189_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__and2_0
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1832_ _1341_ _1335_ net69 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
X_1694_ net21 VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__inv_1
X_1763_ _1106_ _1110_ net68 VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1815_ net30 _1268_ net33 VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1746_ net57 _1064_ net66 VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__mux2_1
X_1677_ _0873_ net114 net68 VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1531_ _0453_ _0451_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__and2_0
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1600_ _0660_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1462_ _0248_ _0246_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__xor2_1
X_1393_ _0051_ _0052_ _0055_ _0058_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_37_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1729_ _0580_ _1033_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__and2_0
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1514_ _0412_ _0410_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__and2_0
X_1445_ _0207_ _0205_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_4_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1428_ net2 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__inv_1
XFILLER_0_33_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1831_ _1324_ net125 net68 VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__mux2_1
X_1621__110 VGND VGND VPWR VPWR _1621__110/HI net110 sky130_fd_sc_hd__conb_1
XFILLER_0_32_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1762_ _1136_ _1130_ net69 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_1
X_1693_ _0901_ _0905_ net68 VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1745_ net24 _1063_ net33 VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__mux2_1
X_1814_ _1236_ _1279_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ net52 _0859_ net66 VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1761__120 VGND VGND VPWR VPWR _1761__120/HI net120 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_14_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1530_ _0455_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1461_ _0248_ _0246_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__and2_0
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1392_ _0032_ _0033_ _0034_ _0035_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_37_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1728_ _1027_ _1025_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1659_ _0785_ _0828_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__and2_0
XFILLER_0_6_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1513_ net41 VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__inv_1
X_1444_ _0207_ _0205_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__and2_0
XFILLER_0_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1537__135 VGND VGND VPWR VPWR _1537__135/HI net135 sky130_fd_sc_hd__conb_1
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1427_ _0122_ _0126_ net68 VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1761_ _1119_ net120 net68 VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux2_1
X_1830_ net64 _1310_ net66 VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1692_ _0931_ _0925_ net69 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1744_ _0990_ _1074_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1813_ _1236_ _1279_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__and2_0
X_1675_ net19 _0858_ net33 VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1391_ _0073_ _0045_ _0047_ _0048_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__nor4_1
X_1460_ _0250_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XTAP_TAPCELL_ROW_37_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1727_ _1027_ _1025_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__and2_0
XFILLER_0_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1658_ _0822_ _0820_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__xor2_1
X_1589_ _0539_ _0623_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__and2_0
XFILLER_0_6_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1512_ net8 VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__inv_1
X_1443_ net36 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__inv_1
XFILLER_0_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1426_ _0152_ _0146_ net69 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1409_ net1 _0079_ net33 VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1760_ net59 _1105_ net66 VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__mux2_1
X_1691_ _0914_ net115 net68 VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1743_ _0990_ _1074_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__and2_0
XFILLER_0_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1674_ _0826_ _0869_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__xor2_1
X_1812_ _1273_ _1271_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_32_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ _0054_ _0065_ _0069_ _0072_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__nor4_1
X_1726_ _1029_ _1030_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1657_ _0822_ _0820_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__and2_0
X_1588_ _0617_ _0615_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1442_ net3 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__inv_1
X_1511_ _0368_ _0372_ net68 VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1709_ net55 VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_0_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1425_ _0108_ net127 net68 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1408_ net67 _0090_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1677__114 VGND VGND VPWR VPWR _1677__114/HI net114 sky130_fd_sc_hd__conb_1
X_1690_ net53 _0900_ net66 VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1811_ _1273_ _1271_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__and2_0
XTAP_TAPCELL_ROW_25_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1742_ _1068_ _1066_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__xor2_1
X_1673_ _0826_ _0869_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__and2_0
XFILLER_0_30_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1725_ _1027_ _1025_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1656_ _0824_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1587_ _0617_ _0615_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__and2_0
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1441_ _0163_ _0167_ net68 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux2_1
X_1510_ _0398_ _0392_ net69 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ net22 VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__inv_1
XFILLER_0_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1639_ net50 VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__inv_1
XFILLER_0_36_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1424_ net58 _0121_ net66 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1407_ net67 _0090_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__and2_0
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1741_ _1068_ _1066_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__and2_0
X_1810_ _1275_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XTAP_TAPCELL_ROW_25_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1672_ _0863_ _0861_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__xor2_1
X_1939_ _0064_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1724_ _1027_ _1025_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__and2_0
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1655_ _0822_ _0820_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1586_ _0619_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_8_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1440_ _0193_ _0187_ net69 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1707_ _0942_ _0946_ net68 VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__mux2_1
X_1638_ net17 VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__inv_1
XFILLER_0_30_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1569_ net45 VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__inv_1
XFILLER_0_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1423_ net25 _0120_ net33 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1406_ _0084_ _0082_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1453__129 VGND VGND VPWR VPWR _1453__129/HI net129 sky130_fd_sc_hd__conb_1
XFILLER_0_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1740_ _1070_ _1071_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1671_ _0863_ _0861_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__and2_0
XFILLER_0_16_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1938_ _0063_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ net56 VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__inv_1
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1654_ _0822_ _0820_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__and2_0
XTAP_TAPCELL_ROW_5_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1585_ _0617_ _0615_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XTAP_TAPCELL_ROW_36_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1706_ _0972_ _0966_ net69 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__mux2_1
X_1637_ _0737_ _0741_ net68 VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__mux2_1
X_1568_ net12 VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__inv_1
X_1499_ net40 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__inv_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1422_ _0030_ _0131_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1495__132 VGND VGND VPWR VPWR _1495__132/HI net132 sky130_fd_sc_hd__conb_1
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1405_ _0084_ _0082_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__and2_0
XFILLER_0_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 a[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1670_ _0865_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1937_ _0062_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1799_ _1195_ _1238_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__and2_0
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ net23 VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__inv_1
XFILLER_0_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1653_ net51 VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__inv_1
X_1584_ _0617_ _0615_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__and2_0
XTAP_TAPCELL_ROW_5_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1705__116 VGND VGND VPWR VPWR _1705__116/HI net116 sky130_fd_sc_hd__conb_1
X_1705_ _0955_ net116 net68 VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1567_ _0532_ _0536_ net68 VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__mux2_1
X_1636_ _0767_ _0761_ net69 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux2_1
X_1498_ net7 VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__inv_1
XFILLER_0_29_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1421_ _0030_ _0131_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__and2_0
XFILLER_0_41_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1619_ net15 _0694_ net33 VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1845__126 VGND VGND VPWR VPWR _1845__126/HI net126 sky130_fd_sc_hd__conb_1
X_1404_ _0086_ _0087_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_23_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 a[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1936_ _0061_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput60 b[4] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
X_1798_ _1232_ _1230_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1721_ _0983_ _0987_ net68 VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593__108 VGND VGND VPWR VPWR _1593__108/HI net108 sky130_fd_sc_hd__conb_1
XFILLER_0_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1652_ net18 VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__inv_1
X_1583_ net46 VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__inv_1
XFILLER_0_21_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1919_ _0074_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1704_ net54 _0941_ net66 VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1566_ _0562_ _0556_ net69 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_1
X_1497_ _0327_ _0331_ net68 VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux2_1
X_1635_ _0750_ net111 net68 VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1420_ _0125_ _0123_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1618_ _0662_ _0705_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__xor2_1
X_1549_ net10 _0489_ net33 VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1403_ _0084_ _0082_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 a[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1935_ _0060_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
Xinput50 b[24] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
Xinput61 b[5] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
X_1797_ _1232_ _1230_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__and2_0
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1720_ _1013_ _1007_ net69 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_1
X_1651_ _0778_ _0782_ net68 VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1582_ net13 VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_36_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1918_ _0073_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1703_ net21 _0940_ net33 VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__mux2_1
X_1634_ net49 _0736_ net66 VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1565_ _0545_ net106 net68 VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__mux2_1
X_1496_ _0357_ _0351_ net69 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1617_ _0662_ _0705_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__and2_0
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1479_ net5 _0284_ net33 VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
X_1548_ _0457_ _0500_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1402_ _0084_ _0082_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__and2_0
XFILLER_0_23_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 a[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1934_ _0059_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput40 b[15] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
X_1796_ _1234_ _1235_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__lpflow_inputiso1p_1
Xinput62 b[6] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
Xinput51 b[25] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1523__134 VGND VGND VPWR VPWR _1523__134/HI net134 sky130_fd_sc_hd__conb_1
X_1581_ _0573_ _0577_ net68 VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__mux2_1
X_1650_ _0808_ _0802_ net69 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1917_ _0072_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_14_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1779_ net61 VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__inv_1
X_1564_ net44 _0531_ net66 VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__mux2_1
X_1702_ _0908_ _0951_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__xor2_1
X_1633_ net16 _0735_ net33 VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1495_ _0340_ net132 net68 VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1547_ _0457_ _0500_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__and2_0
X_1616_ _0699_ _0697_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__xor2_1
X_1478_ _0252_ _0295_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1401_ net34 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_1
XFILLER_0_23_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 a[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1933_ _0058_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput30 a[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
Xinput63 b[7] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
Xinput52 b[26] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
X_1795_ _1232_ _1230_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__lpflow_inputiso1p_1
Xinput41 b[16] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_39_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _0603_ _0597_ net69 VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1916_ _0071_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
X_1847_ _1352_ _1356_ net68 VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1778_ net28 VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_31_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1701_ _0908_ _0951_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__and2_0
XFILLER_0_39_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1494_ net39 _0326_ net66 VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_1
X_1563_ net11 _0530_ net33 VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__mux2_1
X_1632_ _0703_ _0746_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1546_ _0494_ _0492_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__xor2_1
X_1477_ _0252_ _0295_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__and2_0
X_1615_ _0699_ _0697_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__and2_0
XFILLER_0_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1400_ net1 VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_1
Xinput6 a[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_1529_ _0453_ _0451_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput20 a[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_16_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput31 a[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
X_1932_ _0057_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
Xinput42 b[17] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput53 b[27] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
X_1794_ _1232_ _1230_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__and2_0
Xinput64 b[8] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_39_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1777_ _1147_ _1151_ net68 VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1915_ _0070_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
X_1846_ _1382_ _1376_ net69 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1700_ _0945_ _0943_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__xor2_1
X_1631_ _0703_ _0746_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__and2_0
X_1493_ net6 _0325_ net33 VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__mux2_1
X_1562_ _0498_ _0541_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1829_ net31 _1309_ net33 VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__mux2_1
X_1663__113 VGND VGND VPWR VPWR _1663__113/HI net113 sky130_fd_sc_hd__conb_1
XFILLER_0_35_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1614_ _0701_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1476_ _0289_ _0287_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__xor2_1
X_1545_ _0494_ _0492_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and2_0
XFILLER_0_17_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 a[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_1528_ _0453_ _0451_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__and2_0
X_1459_ _0248_ _0246_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1439__128 VGND VGND VPWR VPWR _1439__128/HI net128 sky130_fd_sc_hd__conb_1
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput43 b[18] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput10 a[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput54 b[28] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xinput21 a[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
X_1793_ net62 VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__inv_1
XFILLER_0_24_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput32 a[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
X_1931_ _0056_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
Xinput65 b[9] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1914_ _0069_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
X_1776_ _1177_ _1171_ net69 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1845_ _1365_ net126 net68 VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1630_ _0740_ _0738_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ _0498_ _0541_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__and2_0
X_1492_ _0293_ _0336_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1759_ net26 _1104_ net33 VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__mux2_1
X_1828_ _1277_ _1320_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1544_ _0496_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1613_ _0699_ _0697_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1475_ _0289_ _0287_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__and2_0
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 a[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
X_1527_ net42 VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__inv_1
X_1458_ _0248_ _0246_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__and2_0
X_1389_ _0060_ _0061_ _0063_ _0067_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__nor4_1
XFILLER_0_9_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ _0055_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput33 ainv VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_12
Xinput44 b[19] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput66 binv VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_12
Xinput11 a[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput22 a[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput55 b[29] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1792_ net29 VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__inv_1
XFILLER_0_24_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1913_ _0068_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1775_ _1160_ net121 net68 VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__mux2_1
X_1844_ net65 _1351_ net66 VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1560_ _0535_ _0533_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1491_ _0293_ _0336_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__and2_0
XFILLER_0_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1827_ _1277_ _1320_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__and2_0
XFILLER_0_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1758_ _1031_ _1115_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__xor2_1
X_1689_ net20 _0899_ net33 VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1543_ _0494_ _0492_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1474_ _0291_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1612_ _0699_ _0697_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__and2_0
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 a[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1526_ net9 VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__inv_1
X_1457_ net37 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__inv_1
X_1388_ _0050_ _0053_ _0056_ _0057_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__nor4_1
XFILLER_0_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1509_ _0381_ net133 net68 VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput45 b[1] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput23 a[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput56 b[2] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
Xinput34 b[0] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput12 a[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput67 cin VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_1
X_1791_ _1188_ _1192_ net68 VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__mux2_1
X_1579__107 VGND VGND VPWR VPWR _1579__107/HI net107 sky130_fd_sc_hd__conb_1
XFILLER_0_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1912_ _0065_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
X_1843_ net32 _1350_ net33 VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1774_ net60 _1146_ net66 VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1481__131 VGND VGND VPWR VPWR _1481__131/HI net131 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_41_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1490_ _0330_ _0328_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1826_ _1314_ _1312_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1757_ _1031_ _1115_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__and2_0
X_1688_ _0867_ _0910_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1611_ net48 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__inv_1
XFILLER_0_26_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1473_ _0289_ _0287_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1542_ _0494_ _0492_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__and2_0
XFILLER_0_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1809_ _1273_ _1271_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_31_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1456_ net4 VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__inv_1
X_1525_ _0409_ _0413_ net68 VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput100 net100 VGND VGND VPWR VPWR result[6] sky130_fd_sc_hd__buf_1
X_1508_ net40 _0367_ net66 VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux2_1
X_1439_ _0176_ net128 net68 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput13 a[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
X_1790_ _1218_ _1212_ net69 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_1
Xinput46 b[20] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput68 select[0] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_12
Xinput24 a[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput57 b[30] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput35 b[10] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1911_ _0054_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
X_1773_ net27 _1145_ net33 VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__mux2_1
X_1842_ _1318_ _1361_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_4_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1831__125 VGND VGND VPWR VPWR _1831__125/HI net125 sky130_fd_sc_hd__conb_1
X_1756_ _1109_ _1107_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__xor2_1
X_1825_ _1314_ _1312_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__and2_0
X_1687_ _0867_ _0910_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__and2_0
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1610_ net15 VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__inv_1
XFILLER_0_26_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1541_ net43 VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__inv_1
X_1472_ _0289_ _0287_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__and2_0
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1739_ _1068_ _1066_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1808_ _1273_ _1271_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__and2_0
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1524_ _0439_ _0433_ net69 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux2_1
X_1455_ _0204_ _0208_ net68 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput101 net101 VGND VGND VPWR VPWR result[7] sky130_fd_sc_hd__buf_1
X_1507_ net7 _0366_ net33 VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1438_ net35 _0162_ net66 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput36 b[11] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 a[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 a[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput58 b[31] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xinput47 b[21] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
Xinput69 select[1] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_12
X_1509__133 VGND VGND VPWR VPWR _1509__133/HI net133 sky130_fd_sc_hd__conb_1
XFILLER_0_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1910_ _0043_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1772_ _1113_ _1156_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__xor2_1
X_1841_ _1318_ _1361_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__and2_0
XFILLER_0_34_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1755_ _1109_ _1107_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__and2_0
X_1686_ _0904_ _0902_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1824_ _1316_ _1317_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1540_ net10 VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__inv_1
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1471_ net38 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__inv_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1807_ net63 VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__inv_1
XFILLER_0_32_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1738_ _1068_ _1066_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__and2_0
X_1669_ _0863_ _0861_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1523_ _0422_ net134 net68 VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux2_1
X_1454_ _0234_ _0228_ net69 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput102 net102 VGND VGND VPWR VPWR result[8] sky130_fd_sc_hd__buf_1
XFILLER_0_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1437_ net2 _0161_ net33 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
X_1506_ _0334_ _0377_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput37 b[12] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput26 a[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput59 b[3] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
Xinput48 b[22] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xinput15 a[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_26_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1840_ _1355_ _1353_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1771_ _1113_ _1156_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__and2_0
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1823_ _1314_ _1312_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1754_ _1111_ _1112_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1685_ _0904_ _0902_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__and2_0
XPHY_EDGE_ROW_29_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1470_ net5 VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__inv_1
XFILLER_0_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1806_ net30 VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__inv_1
XFILLER_0_32_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1737_ net57 VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__inv_1
X_1668_ _0863_ _0861_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__and2_0
X_1599_ _0658_ _0656_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1607__109 VGND VGND VPWR VPWR _1607__109/HI net109 sky130_fd_sc_hd__conb_1
X_1522_ net41 _0408_ net66 VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
X_1453_ _0217_ net129 net68 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput103 net103 VGND VGND VPWR VPWR result[9] sky130_fd_sc_hd__buf_1
XFILLER_0_10_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1436_ _0178_ _0172_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__xor2_1
X_1505_ _0334_ _0377_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__and2_0
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1747__119 VGND VGND VPWR VPWR _1747__119/HI net119 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_1_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput38 b[13] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput16 a[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
Xinput27 a[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput49 b[23] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_15_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1419_ _0125_ _0123_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__and2_0
XTAP_TAPCELL_ROW_38_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1770_ _1150_ _1148_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1649__112 VGND VGND VPWR VPWR _1649__112/HI net112 sky130_fd_sc_hd__conb_1
X_1753_ _1109_ _1107_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1822_ _1314_ _1312_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__and2_0
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1684_ _0906_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1736_ net24 VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__inv_1
X_1805_ _1229_ _1233_ net68 VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1667_ net52 VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__inv_1
X_1598_ _0658_ _0656_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__and2_0
XFILLER_0_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1789__122 VGND VGND VPWR VPWR _1789__122/HI net122 sky130_fd_sc_hd__conb_1
XFILLER_0_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1452_ net36 _0203_ net66 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__mux2_1
X_1521_ net8 _0407_ net33 VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1719_ _0996_ net117 net68 VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput104 net104 VGND VGND VPWR VPWR zero sky130_fd_sc_hd__buf_1
XFILLER_0_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1504_ _0371_ _0369_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__xor2_1
X_1435_ _0178_ _0172_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__and2_0
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput39 b[14] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput28 a[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 a[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XFILLER_0_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1418_ _0127_ _0128_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1752_ _1109_ _1107_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__and2_0
X_1683_ _0904_ _0902_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1821_ net64 VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__inv_1
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1735_ _1024_ _1028_ net68 VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__mux2_1
X_1804_ _1259_ _1253_ net69 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_1
X_1666_ net19 VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__inv_1
X_1597_ net47 VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__inv_1
X_1520_ _0375_ _0418_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__xor2_1
X_1451_ net3 _0202_ net33 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1718_ net55 _0982_ net66 VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__mux2_1
X_1649_ _0791_ net112 net68 VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1503_ _0371_ _0369_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__and2_0
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1434_ _0166_ _0164_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_18_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 a[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput29 a[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
XFILLER_0_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1417_ _0125_ _0123_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1820_ net31 VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_32_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1751_ net59 VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__inv_1
X_1682_ _0904_ _0902_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__and2_0
XFILLER_0_24_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1425__127 VGND VGND VPWR VPWR _1425__127/HI net127 sky130_fd_sc_hd__conb_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1803_ _1242_ net123 net68 VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1734_ _1054_ _1048_ net69 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_1
X_1665_ _0819_ _0823_ net68 VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__mux2_1
X_1596_ net14 VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1450_ _0170_ _0213_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__xor2_1
X_1579_ _0586_ net107 net68 VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1717_ net22 _0981_ net33 VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__mux2_1
X_1648_ net50 _0777_ net66 VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1433_ _0166_ _0164_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__and2_0
X_1502_ _0373_ _0374_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XTAP_TAPCELL_ROW_18_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 a[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1416_ _0125_ _0123_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__and2_0
XPHY_EDGE_ROW_5_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1467__130 VGND VGND VPWR VPWR _1467__130/HI net130 sky130_fd_sc_hd__conb_1
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ net26 VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__inv_1
XFILLER_0_29_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1681_ net53 VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__inv_1
XFILLER_0_20_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1733_ _1037_ net118 net68 VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__mux2_1
X_1802_ net62 _1228_ net66 VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1664_ _0849_ _0843_ net69 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__mux2_1
X_1595_ _0614_ _0618_ net68 VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1716_ _0949_ _0992_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1578_ net45 _0572_ net66 VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__mux2_1
X_1647_ net17 _0776_ net33 VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1432_ _0168_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1501_ _0371_ _0369_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XTAP_TAPCELL_ROW_18_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1415_ net58 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1817__124 VGND VGND VPWR VPWR _1817__124/HI net124 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1680_ net20 VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__inv_1
XFILLER_0_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1732_ net56 _1023_ net66 VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__mux2_1
X_1663_ _0832_ net113 net68 VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__mux2_1
X_1801_ net29 _1227_ net33 VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1594_ _0644_ _0638_ net69 VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1715_ _0949_ _0992_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__and2_0
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1646_ _0744_ _0787_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__xor2_1
X_1565__106 VGND VGND VPWR VPWR _1565__106/HI net106 sky130_fd_sc_hd__conb_1
XFILLER_0_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1577_ net12 _0571_ net33 VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1500_ _0371_ _0369_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__and2_0
Xoutput90 net90 VGND VGND VPWR VPWR result[26] sky130_fd_sc_hd__buf_1
X_1431_ _0166_ _0164_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XTAP_TAPCELL_ROW_18_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1629_ _0740_ _0738_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__and2_0
XFILLER_0_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1414_ net25 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_6_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1800_ _1195_ _1238_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1731_ net23 _1022_ net33 VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__mux2_1
X_1662_ net51 _0818_ net66 VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1593_ _0627_ net108 net68 VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1929_ _0053_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1576_ _0088_ _0582_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__xor2_1
X_1714_ _0986_ _0984_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1645_ _0744_ _0787_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__and2_0
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1430_ _0166_ _0164_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__and2_0
Xoutput80 net80 VGND VGND VPWR VPWR result[17] sky130_fd_sc_hd__buf_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput91 net91 VGND VGND VPWR VPWR result[27] sky130_fd_sc_hd__buf_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1559_ _0535_ _0533_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__and2_0
XFILLER_0_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1628_ _0742_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1413_ _0081_ _0085_ net68 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1730_ _0580_ _1033_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1661_ net18 _0817_ net33 VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1592_ net46 _0613_ net66 VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1928_ _0052_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1713_ _0986_ _0984_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__and2_0
X_1575_ _0088_ _0582_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__and2_0
X_1644_ _0781_ _0779_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput70 net70 VGND VGND VPWR VPWR cout sky130_fd_sc_hd__buf_1
XFILLER_0_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput81 net81 VGND VGND VPWR VPWR result[18] sky130_fd_sc_hd__buf_1
XFILLER_0_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput92 net92 VGND VGND VPWR VPWR result[28] sky130_fd_sc_hd__buf_1
XFILLER_0_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1558_ _0537_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1489_ _0330_ _0328_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__and2_0
X_1627_ _0740_ _0738_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1412_ _0111_ _0105_ net69 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1660_ _0785_ _0828_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__xor2_1
X_1591_ net13 _0612_ net33 VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1927_ _0051_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
X_1789_ _1201_ net122 net68 VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__mux2_1
X_1712_ _0988_ _0989_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1643_ _0781_ _0779_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__and2_0
X_1574_ _0576_ _0574_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput93 net93 VGND VGND VPWR VPWR result[29] sky130_fd_sc_hd__buf_1
Xoutput71 net71 VGND VGND VPWR VPWR overflow sky130_fd_sc_hd__buf_1
Xoutput82 net82 VGND VGND VPWR VPWR result[19] sky130_fd_sc_hd__buf_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1626_ _0740_ _0738_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__and2_0
X_1557_ _0535_ _0533_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1488_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1411_ _0094_ _0108_ net68 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1609_ _0655_ _0659_ net68 VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ _0539_ _0623_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__xor2_1
X_1788_ net61 _1187_ net66 VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1926_ _0050_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
X_1733__118 VGND VGND VPWR VPWR _1733__118/HI net118 sky130_fd_sc_hd__conb_1
XFILLER_0_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1711_ _0986_ _0984_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1642_ _0783_ _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1573_ _0576_ _0574_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__and2_0
XFILLER_0_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput94 net94 VGND VGND VPWR VPWR result[2] sky130_fd_sc_hd__buf_1
Xoutput83 net83 VGND VGND VPWR VPWR result[1] sky130_fd_sc_hd__buf_1
Xoutput72 net72 VGND VGND VPWR VPWR result[0] sky130_fd_sc_hd__buf_1
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1556_ _0535_ _0533_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__and2_0
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1625_ net49 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__inv_1
X_1487_ _0330_ _0328_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__lpflow_inputiso1p_1
XFILLER_0_27_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1410_ net34 _0080_ net66 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1635__111 VGND VGND VPWR VPWR _1635__111/HI net111 sky130_fd_sc_hd__conb_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1539_ _0450_ _0454_ net68 VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux2_1
X_1608_ _0685_ _0679_ net69 VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1775__121 VGND VGND VPWR VPWR _1775__121/HI net121 sky130_fd_sc_hd__conb_1
XFILLER_0_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1925_ _0049_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
X_1787_ net28 _1186_ net33 VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1572_ _0578_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1710_ _0986_ _0984_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__and2_0
XFILLER_0_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1641_ _0781_ _0779_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1839_ _1355_ _1353_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__and2_0
XFILLER_0_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput95 net95 VGND VGND VPWR VPWR result[30] sky130_fd_sc_hd__buf_1
Xoutput73 net73 VGND VGND VPWR VPWR result[10] sky130_fd_sc_hd__buf_1
Xoutput84 net84 VGND VGND VPWR VPWR result[20] sky130_fd_sc_hd__buf_1
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1555_ net44 VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__inv_1
X_1624_ net16 VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__inv_1
X_1486_ _0330_ _0328_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__and2_0
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1538_ _0480_ _0474_ net69 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1607_ _0668_ net109 net68 VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux2_1
X_1469_ _0245_ _0249_ net68 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1941_ _0067_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1924_ _0048_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
X_1786_ _1154_ _1197_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1571_ _0576_ _0574_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1640_ _0781_ _0779_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__and2_0
XFILLER_0_21_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1838_ _1357_ _1358_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__lpflow_inputiso1p_1
X_1769_ _1150_ _1148_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__and2_0
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput74 net74 VGND VGND VPWR VPWR result[11] sky130_fd_sc_hd__buf_1
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput96 net96 VGND VGND VPWR VPWR result[31] sky130_fd_sc_hd__buf_1
Xoutput85 net85 VGND VGND VPWR VPWR result[21] sky130_fd_sc_hd__buf_1
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1485_ net39 VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__inv_1
X_1554_ net11 VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__inv_1
X_1623_ _0696_ _0700_ net68 VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__mux2_1
.ends

