magic
tech sky130A
magscale 1 2
timestamp 1743984716
<< nwell >>
rect 1066 2159 24050 25041
<< obsli1 >>
rect 1104 2159 24012 25041
<< obsm1 >>
rect 842 2128 24072 25072
<< metal2 >>
rect 5814 26516 5870 27316
rect 6458 26516 6514 27316
rect 7102 26516 7158 27316
rect 7746 26516 7802 27316
rect 8390 26516 8446 27316
rect 9034 26516 9090 27316
rect 9678 26516 9734 27316
rect 10322 26516 10378 27316
rect 10966 26516 11022 27316
rect 11610 26516 11666 27316
rect 12254 26516 12310 27316
rect 12898 26516 12954 27316
rect 13542 26516 13598 27316
rect 14186 26516 14242 27316
rect 14830 26516 14886 27316
rect 15474 26516 15530 27316
rect 16118 26516 16174 27316
rect 16762 26516 16818 27316
rect 17406 26516 17462 27316
rect 18050 26516 18106 27316
rect 20626 26516 20682 27316
rect 18 0 74 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
<< obsm2 >>
rect 846 26460 5758 26602
rect 5926 26460 6402 26602
rect 6570 26460 7046 26602
rect 7214 26460 7690 26602
rect 7858 26460 8334 26602
rect 8502 26460 8978 26602
rect 9146 26460 9622 26602
rect 9790 26460 10266 26602
rect 10434 26460 10910 26602
rect 11078 26460 11554 26602
rect 11722 26460 12198 26602
rect 12366 26460 12842 26602
rect 13010 26460 13486 26602
rect 13654 26460 14130 26602
rect 14298 26460 14774 26602
rect 14942 26460 15418 26602
rect 15586 26460 16062 26602
rect 16230 26460 16706 26602
rect 16874 26460 17350 26602
rect 17518 26460 17994 26602
rect 18162 26460 20570 26602
rect 20738 26460 23900 26602
rect 846 856 23900 26460
rect 846 734 3182 856
rect 3350 734 3826 856
rect 3994 734 4470 856
rect 4638 734 5114 856
rect 5282 734 5758 856
rect 5926 734 6402 856
rect 6570 734 7046 856
rect 7214 734 7690 856
rect 7858 734 8334 856
rect 8502 734 8978 856
rect 9146 734 9622 856
rect 9790 734 10266 856
rect 10434 734 10910 856
rect 11078 734 11554 856
rect 11722 734 12198 856
rect 12366 734 12842 856
rect 13010 734 13486 856
rect 13654 734 14130 856
rect 14298 734 14774 856
rect 14942 734 15418 856
rect 15586 734 16062 856
rect 16230 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17994 856
rect 18162 734 18638 856
rect 18806 734 19282 856
rect 19450 734 19926 856
rect 20094 734 20570 856
rect 20738 734 21214 856
rect 21382 734 23900 856
<< metal3 >>
rect 24372 24488 25172 24608
rect 24372 23808 25172 23928
rect 24372 23128 25172 23248
rect 24372 22448 25172 22568
rect 24372 21768 25172 21888
rect 0 21088 800 21208
rect 24372 21088 25172 21208
rect 0 20408 800 20528
rect 24372 20408 25172 20528
rect 0 19728 800 19848
rect 24372 19728 25172 19848
rect 0 19048 800 19168
rect 24372 19048 25172 19168
rect 0 18368 800 18488
rect 24372 18368 25172 18488
rect 0 17688 800 17808
rect 24372 17688 25172 17808
rect 0 17008 800 17128
rect 24372 17008 25172 17128
rect 0 16328 800 16448
rect 24372 16328 25172 16448
rect 0 15648 800 15768
rect 24372 15648 25172 15768
rect 0 14968 800 15088
rect 24372 14968 25172 15088
rect 0 14288 800 14408
rect 24372 14288 25172 14408
rect 0 13608 800 13728
rect 24372 13608 25172 13728
rect 0 12928 800 13048
rect 24372 12928 25172 13048
rect 0 12248 800 12368
rect 24372 12248 25172 12368
rect 0 11568 800 11688
rect 24372 11568 25172 11688
rect 0 10888 800 11008
rect 24372 10888 25172 11008
rect 0 10208 800 10328
rect 24372 10208 25172 10328
rect 0 9528 800 9648
rect 24372 9528 25172 9648
rect 0 8848 800 8968
rect 24372 8848 25172 8968
rect 24372 8168 25172 8288
rect 0 7488 800 7608
rect 24372 7488 25172 7608
rect 0 6808 800 6928
rect 24372 6808 25172 6928
rect 24372 6128 25172 6248
rect 24372 5448 25172 5568
rect 24372 4768 25172 4888
rect 24372 4088 25172 4208
rect 24372 3408 25172 3528
rect 24372 2728 25172 2848
<< obsm3 >>
rect 798 24688 24372 25057
rect 798 24408 24292 24688
rect 798 24008 24372 24408
rect 798 23728 24292 24008
rect 798 23328 24372 23728
rect 798 23048 24292 23328
rect 798 22648 24372 23048
rect 798 22368 24292 22648
rect 798 21968 24372 22368
rect 798 21688 24292 21968
rect 798 21288 24372 21688
rect 880 21008 24292 21288
rect 798 20608 24372 21008
rect 880 20328 24292 20608
rect 798 19928 24372 20328
rect 880 19648 24292 19928
rect 798 19248 24372 19648
rect 880 18968 24292 19248
rect 798 18568 24372 18968
rect 880 18288 24292 18568
rect 798 17888 24372 18288
rect 880 17608 24292 17888
rect 798 17208 24372 17608
rect 880 16928 24292 17208
rect 798 16528 24372 16928
rect 880 16248 24292 16528
rect 798 15848 24372 16248
rect 880 15568 24292 15848
rect 798 15168 24372 15568
rect 880 14888 24292 15168
rect 798 14488 24372 14888
rect 880 14208 24292 14488
rect 798 13808 24372 14208
rect 880 13528 24292 13808
rect 798 13128 24372 13528
rect 880 12848 24292 13128
rect 798 12448 24372 12848
rect 880 12168 24292 12448
rect 798 11768 24372 12168
rect 880 11488 24292 11768
rect 798 11088 24372 11488
rect 880 10808 24292 11088
rect 798 10408 24372 10808
rect 880 10128 24292 10408
rect 798 9728 24372 10128
rect 880 9448 24292 9728
rect 798 9048 24372 9448
rect 880 8768 24292 9048
rect 798 8368 24372 8768
rect 798 8088 24292 8368
rect 798 7688 24372 8088
rect 880 7408 24292 7688
rect 798 7008 24372 7408
rect 880 6728 24292 7008
rect 798 6328 24372 6728
rect 798 6048 24292 6328
rect 798 5648 24372 6048
rect 798 5368 24292 5648
rect 798 4968 24372 5368
rect 798 4688 24292 4968
rect 798 4288 24372 4688
rect 798 4008 24292 4288
rect 798 3608 24372 4008
rect 798 3328 24292 3608
rect 798 2928 24372 3328
rect 798 2648 24292 2928
rect 798 2143 24372 2648
<< metal4 >>
rect 3807 2128 4127 25072
rect 4467 2128 4787 25072
rect 9534 2128 9854 25072
rect 10194 2128 10514 25072
rect 15261 2128 15581 25072
rect 15921 2128 16241 25072
rect 20988 2128 21308 25072
rect 21648 2128 21968 25072
<< metal5 >>
rect 1056 22668 24060 22988
rect 1056 22008 24060 22328
rect 1056 16956 24060 17276
rect 1056 16296 24060 16616
rect 1056 11244 24060 11564
rect 1056 10584 24060 10904
rect 1056 5532 24060 5852
rect 1056 4872 24060 5192
<< labels >>
rlabel metal4 s 4467 2128 4787 25072 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 10194 2128 10514 25072 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 15921 2128 16241 25072 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 21648 2128 21968 25072 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5532 24060 5852 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 11244 24060 11564 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 16956 24060 17276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 22668 24060 22988 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3807 2128 4127 25072 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9534 2128 9854 25072 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 15261 2128 15581 25072 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 20988 2128 21308 25072 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4872 24060 5192 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 10584 24060 10904 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 16296 24060 16616 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 22008 24060 22328 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 3238 0 3294 800 6 a[0]
port 3 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 a[10]
port 4 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 a[11]
port 5 nsew signal input
rlabel metal2 s 5814 26516 5870 27316 6 a[12]
port 6 nsew signal input
rlabel metal2 s 7746 26516 7802 27316 6 a[13]
port 7 nsew signal input
rlabel metal2 s 12254 26516 12310 27316 6 a[14]
port 8 nsew signal input
rlabel metal2 s 12898 26516 12954 27316 6 a[15]
port 9 nsew signal input
rlabel metal3 s 24372 23128 25172 23248 6 a[16]
port 10 nsew signal input
rlabel metal2 s 16762 26516 16818 27316 6 a[17]
port 11 nsew signal input
rlabel metal2 s 18050 26516 18106 27316 6 a[18]
port 12 nsew signal input
rlabel metal3 s 24372 22448 25172 22568 6 a[19]
port 13 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 a[1]
port 14 nsew signal input
rlabel metal3 s 24372 21768 25172 21888 6 a[20]
port 15 nsew signal input
rlabel metal3 s 24372 16328 25172 16448 6 a[21]
port 16 nsew signal input
rlabel metal3 s 24372 14968 25172 15088 6 a[22]
port 17 nsew signal input
rlabel metal3 s 24372 4768 25172 4888 6 a[23]
port 18 nsew signal input
rlabel metal3 s 24372 11568 25172 11688 6 a[24]
port 19 nsew signal input
rlabel metal3 s 24372 12248 25172 12368 6 a[25]
port 20 nsew signal input
rlabel metal3 s 24372 5448 25172 5568 6 a[26]
port 21 nsew signal input
rlabel metal3 s 24372 6128 25172 6248 6 a[27]
port 22 nsew signal input
rlabel metal3 s 24372 2728 25172 2848 6 a[28]
port 23 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 a[29]
port 24 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 a[2]
port 25 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 a[30]
port 26 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 a[31]
port 27 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 a[3]
port 28 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 a[4]
port 29 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 a[5]
port 30 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 a[6]
port 31 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 a[7]
port 32 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 a[8]
port 33 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 a[9]
port 34 nsew signal input
rlabel metal3 s 24372 24488 25172 24608 6 ainv
port 35 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 b[0]
port 36 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 b[10]
port 37 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 b[11]
port 38 nsew signal input
rlabel metal2 s 6458 26516 6514 27316 6 b[12]
port 39 nsew signal input
rlabel metal2 s 7102 26516 7158 27316 6 b[13]
port 40 nsew signal input
rlabel metal2 s 11610 26516 11666 27316 6 b[14]
port 41 nsew signal input
rlabel metal2 s 13542 26516 13598 27316 6 b[15]
port 42 nsew signal input
rlabel metal3 s 24372 18368 25172 18488 6 b[16]
port 43 nsew signal input
rlabel metal2 s 14830 26516 14886 27316 6 b[17]
port 44 nsew signal input
rlabel metal2 s 17406 26516 17462 27316 6 b[18]
port 45 nsew signal input
rlabel metal2 s 20626 26516 20682 27316 6 b[19]
port 46 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 b[1]
port 47 nsew signal input
rlabel metal3 s 24372 20408 25172 20528 6 b[20]
port 48 nsew signal input
rlabel metal3 s 24372 15648 25172 15768 6 b[21]
port 49 nsew signal input
rlabel metal3 s 24372 14288 25172 14408 6 b[22]
port 50 nsew signal input
rlabel metal3 s 24372 13608 25172 13728 6 b[23]
port 51 nsew signal input
rlabel metal3 s 24372 10888 25172 11008 6 b[24]
port 52 nsew signal input
rlabel metal3 s 24372 12928 25172 13048 6 b[25]
port 53 nsew signal input
rlabel metal3 s 24372 10208 25172 10328 6 b[26]
port 54 nsew signal input
rlabel metal3 s 24372 7488 25172 7608 6 b[27]
port 55 nsew signal input
rlabel metal3 s 24372 3408 25172 3528 6 b[28]
port 56 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 b[29]
port 57 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 b[2]
port 58 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 b[30]
port 59 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 b[31]
port 60 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 b[3]
port 61 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 b[4]
port 62 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 b[5]
port 63 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 b[6]
port 64 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 b[7]
port 65 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 b[8]
port 66 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 b[9]
port 67 nsew signal input
rlabel metal3 s 24372 23808 25172 23928 6 binv
port 68 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 cin
port 69 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 cout
port 70 nsew signal output
rlabel metal2 s 18 0 74 800 6 fake_clk
port 71 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 overflow
port 72 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 result[0]
port 73 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 result[10]
port 74 nsew signal output
rlabel metal2 s 8390 26516 8446 27316 6 result[11]
port 75 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 result[12]
port 76 nsew signal output
rlabel metal2 s 9034 26516 9090 27316 6 result[13]
port 77 nsew signal output
rlabel metal2 s 10322 26516 10378 27316 6 result[14]
port 78 nsew signal output
rlabel metal2 s 9678 26516 9734 27316 6 result[15]
port 79 nsew signal output
rlabel metal3 s 24372 17688 25172 17808 6 result[16]
port 80 nsew signal output
rlabel metal2 s 14186 26516 14242 27316 6 result[17]
port 81 nsew signal output
rlabel metal2 s 16118 26516 16174 27316 6 result[18]
port 82 nsew signal output
rlabel metal3 s 24372 19728 25172 19848 6 result[19]
port 83 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 result[1]
port 84 nsew signal output
rlabel metal3 s 24372 19048 25172 19168 6 result[20]
port 85 nsew signal output
rlabel metal3 s 24372 17008 25172 17128 6 result[21]
port 86 nsew signal output
rlabel metal3 s 24372 21088 25172 21208 6 result[22]
port 87 nsew signal output
rlabel metal2 s 15474 26516 15530 27316 6 result[23]
port 88 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 result[24]
port 89 nsew signal output
rlabel metal3 s 24372 6808 25172 6928 6 result[25]
port 90 nsew signal output
rlabel metal3 s 24372 9528 25172 9648 6 result[26]
port 91 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 result[27]
port 92 nsew signal output
rlabel metal3 s 24372 8848 25172 8968 6 result[28]
port 93 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 result[29]
port 94 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 result[2]
port 95 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 result[30]
port 96 nsew signal output
rlabel metal3 s 24372 8168 25172 8288 6 result[31]
port 97 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 result[3]
port 98 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 result[4]
port 99 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 result[5]
port 100 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 result[6]
port 101 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 result[7]
port 102 nsew signal output
rlabel metal2 s 10966 26516 11022 27316 6 result[8]
port 103 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 result[9]
port 104 nsew signal output
rlabel metal3 s 24372 4088 25172 4208 6 select[0]
port 105 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 select[1]
port 106 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 zero
port 107 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 25172 27316
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1364238
string GDS_FILE /home/prajuval/Desktop/OpenLane/openlane/n_bit_alu/runs/run_11/results/signoff/n_bit_alu.magic.gds
string GDS_START 81026
<< end >>

